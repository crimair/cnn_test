// soc_system_mem_0.v

// Generated using ACDS version 13.1 162 at 2015.04.08.02:28:25

`timescale 1 ps / 1 ps
module soc_system_mem_0 (
		input  wire         clk_clk,                                                  //                            clk.clk
		input  wire         reset_reset_n,                                            //                          reset.reset_n
		output wire [14:0]  memory_0_mem_a,                                           //                       memory_0.mem_a
		output wire [2:0]   memory_0_mem_ba,                                          //                               .mem_ba
		output wire [0:0]   memory_0_mem_ck,                                          //                               .mem_ck
		output wire [0:0]   memory_0_mem_ck_n,                                        //                               .mem_ck_n
		output wire [0:0]   memory_0_mem_cke,                                         //                               .mem_cke
		output wire [0:0]   memory_0_mem_cs_n,                                        //                               .mem_cs_n
		output wire [3:0]   memory_0_mem_dm,                                          //                               .mem_dm
		output wire [0:0]   memory_0_mem_ras_n,                                       //                               .mem_ras_n
		output wire [0:0]   memory_0_mem_cas_n,                                       //                               .mem_cas_n
		output wire [0:0]   memory_0_mem_we_n,                                        //                               .mem_we_n
		output wire         memory_0_mem_reset_n,                                     //                               .mem_reset_n
		inout  wire [31:0]  memory_0_mem_dq,                                          //                               .mem_dq
		inout  wire [3:0]   memory_0_mem_dqs,                                         //                               .mem_dqs
		inout  wire [3:0]   memory_0_mem_dqs_n,                                       //                               .mem_dqs_n
		output wire [0:0]   memory_0_mem_odt,                                         //                               .mem_odt
		input  wire         oct_rzqin,                                                //                            oct.rzqin
		output wire         mem_if_ddr3_emif_0_status_local_init_done,                //      mem_if_ddr3_emif_0_status.local_init_done
		output wire         mem_if_ddr3_emif_0_status_local_cal_success,              //                               .local_cal_success
		output wire         mem_if_ddr3_emif_0_status_local_cal_fail,                 //                               .local_cal_fail
		output wire         mem_if_ddr3_emif_0_pll_sharing_pll_mem_clk,               // mem_if_ddr3_emif_0_pll_sharing.pll_mem_clk
		output wire         mem_if_ddr3_emif_0_pll_sharing_pll_write_clk,             //                               .pll_write_clk
		output wire         mem_if_ddr3_emif_0_pll_sharing_pll_locked,                //                               .pll_locked
		output wire         mem_if_ddr3_emif_0_pll_sharing_pll_write_clk_pre_phy_clk, //                               .pll_write_clk_pre_phy_clk
		output wire         mem_if_ddr3_emif_0_pll_sharing_pll_addr_cmd_clk,          //                               .pll_addr_cmd_clk
		output wire         mem_if_ddr3_emif_0_pll_sharing_pll_avl_clk,               //                               .pll_avl_clk
		output wire         mem_if_ddr3_emif_0_pll_sharing_pll_config_clk,            //                               .pll_config_clk
		output wire         mem_if_ddr3_emif_0_pll_sharing_pll_dr_clk,                //                               .pll_dr_clk
		output wire         mem_if_ddr3_emif_0_pll_sharing_pll_dr_clk_pre_phy_clk,    //                               .pll_dr_clk_pre_phy_clk
		output wire         mem_if_ddr3_emif_0_pll_sharing_pll_mem_phy_clk,           //                               .pll_mem_phy_clk
		output wire         mem_if_ddr3_emif_0_pll_sharing_afi_phy_clk,               //                               .afi_phy_clk
		output wire         mem_if_ddr3_emif_0_pll_sharing_pll_avl_phy_clk,           //                               .pll_avl_phy_clk
		output wire         afi_clk_clk,                                              //                        afi_clk.clk
		output wire         mem0_waitrequest,                                         //                           mem0.waitrequest
		output wire [127:0] mem0_readdata,                                            //                               .readdata
		output wire         mem0_readdatavalid,                                       //                               .readdatavalid
		input  wire [2:0]   mem0_burstcount,                                          //                               .burstcount
		input  wire [127:0] mem0_writedata,                                           //                               .writedata
		input  wire [25:0]  mem0_address,                                             //                               .address
		input  wire         mem0_write,                                               //                               .write
		input  wire         mem0_read,                                                //                               .read
		input  wire [15:0]  mem0_byteenable,                                          //                               .byteenable
		input  wire         mem0_debugaccess,                                         //                               .debugaccess
		output wire         mem1_waitrequest,                                         //                           mem1.waitrequest
		output wire [127:0] mem1_readdata,                                            //                               .readdata
		output wire         mem1_readdatavalid,                                       //                               .readdatavalid
		input  wire [2:0]   mem1_burstcount,                                          //                               .burstcount
		input  wire [127:0] mem1_writedata,                                           //                               .writedata
		input  wire [25:0]  mem1_address,                                             //                               .address
		input  wire         mem1_write,                                               //                               .write
		input  wire         mem1_read,                                                //                               .read
		input  wire [15:0]  mem1_byteenable,                                          //                               .byteenable
		input  wire         mem1_debugaccess,                                         //                               .debugaccess
		output wire         mem2_waitrequest,                                         //                           mem2.waitrequest
		output wire [127:0] mem2_readdata,                                            //                               .readdata
		output wire         mem2_readdatavalid,                                       //                               .readdatavalid
		input  wire [2:0]   mem2_burstcount,                                          //                               .burstcount
		input  wire [127:0] mem2_writedata,                                           //                               .writedata
		input  wire [25:0]  mem2_address,                                             //                               .address
		input  wire         mem2_write,                                               //                               .write
		input  wire         mem2_read,                                                //                               .read
		input  wire [15:0]  mem2_byteenable,                                          //                               .byteenable
		input  wire         mem2_debugaccess,                                         //                               .debugaccess
		output wire         mem3_waitrequest,                                         //                           mem3.waitrequest
		output wire [127:0] mem3_readdata,                                            //                               .readdata
		output wire         mem3_readdatavalid,                                       //                               .readdatavalid
		input  wire [2:0]   mem3_burstcount,                                          //                               .burstcount
		input  wire [127:0] mem3_writedata,                                           //                               .writedata
		input  wire [25:0]  mem3_address,                                             //                               .address
		input  wire         mem3_write,                                               //                               .write
		input  wire         mem3_read,                                                //                               .read
		input  wire [15:0]  mem3_byteenable,                                          //                               .byteenable
		input  wire         mem3_debugaccess,                                         //                               .debugaccess
		output wire         mem4_waitrequest,                                         //                           mem4.waitrequest
		output wire [127:0] mem4_readdata,                                            //                               .readdata
		output wire         mem4_readdatavalid,                                       //                               .readdatavalid
		input  wire [2:0]   mem4_burstcount,                                          //                               .burstcount
		input  wire [127:0] mem4_writedata,                                           //                               .writedata
		input  wire [25:0]  mem4_address,                                             //                               .address
		input  wire         mem4_write,                                               //                               .write
		input  wire         mem4_read,                                                //                               .read
		input  wire [15:0]  mem4_byteenable,                                          //                               .byteenable
		input  wire         mem4_debugaccess,                                         //                               .debugaccess
		output wire         cam0_waitrequest,                                         //                           cam0.waitrequest
		output wire [127:0] cam0_readdata,                                            //                               .readdata
		output wire         cam0_readdatavalid,                                       //                               .readdatavalid
		input  wire [2:0]   cam0_burstcount,                                          //                               .burstcount
		input  wire [127:0] cam0_writedata,                                           //                               .writedata
		input  wire [25:0]  cam0_address,                                             //                               .address
		input  wire         cam0_write,                                               //                               .write
		input  wire         cam0_read,                                                //                               .read
		input  wire [15:0]  cam0_byteenable,                                          //                               .byteenable
		input  wire         cam0_debugaccess,                                         //                               .debugaccess
		output wire         cam1_waitrequest,                                         //                           cam1.waitrequest
		output wire [127:0] cam1_readdata,                                            //                               .readdata
		output wire         cam1_readdatavalid,                                       //                               .readdatavalid
		input  wire [2:0]   cam1_burstcount,                                          //                               .burstcount
		input  wire [127:0] cam1_writedata,                                           //                               .writedata
		input  wire [25:0]  cam1_address,                                             //                               .address
		input  wire         cam1_write,                                               //                               .write
		input  wire         cam1_read,                                                //                               .read
		input  wire [15:0]  cam1_byteenable,                                          //                               .byteenable
		input  wire         cam1_debugaccess,                                         //                               .debugaccess
		output wire         cam23_waitrequest,                                        //                          cam23.waitrequest
		output wire [127:0] cam23_readdata,                                           //                               .readdata
		output wire         cam23_readdatavalid,                                      //                               .readdatavalid
		input  wire [2:0]   cam23_burstcount,                                         //                               .burstcount
		input  wire [127:0] cam23_writedata,                                          //                               .writedata
		input  wire [25:0]  cam23_address,                                            //                               .address
		input  wire         cam23_write,                                              //                               .write
		input  wire         cam23_read,                                               //                               .read
		input  wire [15:0]  cam23_byteenable,                                         //                               .byteenable
		input  wire         cam23_debugaccess,                                        //                               .debugaccess
		output wire         cam45_waitrequest,                                        //                          cam45.waitrequest
		output wire [127:0] cam45_readdata,                                           //                               .readdata
		output wire         cam45_readdatavalid,                                      //                               .readdatavalid
		input  wire [2:0]   cam45_burstcount,                                         //                               .burstcount
		input  wire [127:0] cam45_writedata,                                          //                               .writedata
		input  wire [25:0]  cam45_address,                                            //                               .address
		input  wire         cam45_write,                                              //                               .write
		input  wire         cam45_read,                                               //                               .read
		input  wire [15:0]  cam45_byteenable,                                         //                               .byteenable
		input  wire         cam45_debugaccess,                                        //                               .debugaccess
		output wire         hps_waitrequest,                                          //                            hps.waitrequest
		output wire [127:0] hps_readdata,                                             //                               .readdata
		output wire         hps_readdatavalid,                                        //                               .readdatavalid
		input  wire [2:0]   hps_burstcount,                                           //                               .burstcount
		input  wire [127:0] hps_writedata,                                            //                               .writedata
		input  wire [25:0]  hps_address,                                              //                               .address
		input  wire         hps_write,                                                //                               .write
		input  wire         hps_read,                                                 //                               .read
		input  wire [15:0]  hps_byteenable,                                           //                               .byteenable
		input  wire         hps_debugaccess,                                          //                               .debugaccess
		output wire         test_vga_waitrequest,                                     //                       test_vga.waitrequest
		output wire [127:0] test_vga_readdata,                                        //                               .readdata
		output wire         test_vga_readdatavalid,                                   //                               .readdatavalid
		input  wire [2:0]   test_vga_burstcount,                                      //                               .burstcount
		input  wire [127:0] test_vga_writedata,                                       //                               .writedata
		input  wire [25:0]  test_vga_address,                                         //                               .address
		input  wire         test_vga_write,                                           //                               .write
		input  wire         test_vga_read,                                            //                               .read
		input  wire [15:0]  test_vga_byteenable,                                      //                               .byteenable
		input  wire         test_vga_debugaccess,                                     //                               .debugaccess
		input  wire         clk_0_clk                                                 //                          clk_0.clk
	);

	wire          mem_if_ddr3_emif_0_afi_clk_clk;                                // mem_if_ddr3_emif_0:afi_clk -> [mem_if_ddr3_emif_0:mp_cmd_clk_0_clk, mem_if_ddr3_emif_0:mp_rfifo_clk_0_clk, mem_if_ddr3_emif_0:mp_wfifo_clk_0_clk, mm_interconnect_0:mem_if_ddr3_emif_0_afi_clk_clk, rst_controller_002:clk]
	wire          mm_interconnect_0_mem_if_ddr3_emif_0_avl_0_waitrequest;        // mem_if_ddr3_emif_0:avl_ready_0 -> mm_interconnect_0:mem_if_ddr3_emif_0_avl_0_waitrequest
	wire    [1:0] mm_interconnect_0_mem_if_ddr3_emif_0_avl_0_burstcount;         // mm_interconnect_0:mem_if_ddr3_emif_0_avl_0_burstcount -> mem_if_ddr3_emif_0:avl_size_0
	wire   [31:0] mm_interconnect_0_mem_if_ddr3_emif_0_avl_0_writedata;          // mm_interconnect_0:mem_if_ddr3_emif_0_avl_0_writedata -> mem_if_ddr3_emif_0:avl_wdata_0
	wire   [27:0] mm_interconnect_0_mem_if_ddr3_emif_0_avl_0_address;            // mm_interconnect_0:mem_if_ddr3_emif_0_avl_0_address -> mem_if_ddr3_emif_0:avl_addr_0
	wire          mm_interconnect_0_mem_if_ddr3_emif_0_avl_0_write;              // mm_interconnect_0:mem_if_ddr3_emif_0_avl_0_write -> mem_if_ddr3_emif_0:avl_write_req_0
	wire          mm_interconnect_0_mem_if_ddr3_emif_0_avl_0_beginbursttransfer; // mm_interconnect_0:mem_if_ddr3_emif_0_avl_0_beginbursttransfer -> mem_if_ddr3_emif_0:avl_burstbegin_0
	wire          mm_interconnect_0_mem_if_ddr3_emif_0_avl_0_read;               // mm_interconnect_0:mem_if_ddr3_emif_0_avl_0_read -> mem_if_ddr3_emif_0:avl_read_req_0
	wire   [31:0] mm_interconnect_0_mem_if_ddr3_emif_0_avl_0_readdata;           // mem_if_ddr3_emif_0:avl_rdata_0 -> mm_interconnect_0:mem_if_ddr3_emif_0_avl_0_readdata
	wire          mm_interconnect_0_mem_if_ddr3_emif_0_avl_0_readdatavalid;      // mem_if_ddr3_emif_0:avl_rdata_valid_0 -> mm_interconnect_0:mem_if_ddr3_emif_0_avl_0_readdatavalid
	wire    [3:0] mm_interconnect_0_mem_if_ddr3_emif_0_avl_0_byteenable;         // mm_interconnect_0:mem_if_ddr3_emif_0_avl_0_byteenable -> mem_if_ddr3_emif_0:avl_be_0
	wire    [2:0] mm_bridge_9_m0_burstcount;                                     // mm_bridge_9:m0_burstcount -> mm_interconnect_0:mm_bridge_9_m0_burstcount
	wire          mm_bridge_9_m0_waitrequest;                                    // mm_interconnect_0:mm_bridge_9_m0_waitrequest -> mm_bridge_9:m0_waitrequest
	wire   [25:0] mm_bridge_9_m0_address;                                        // mm_bridge_9:m0_address -> mm_interconnect_0:mm_bridge_9_m0_address
	wire  [127:0] mm_bridge_9_m0_writedata;                                      // mm_bridge_9:m0_writedata -> mm_interconnect_0:mm_bridge_9_m0_writedata
	wire          mm_bridge_9_m0_write;                                          // mm_bridge_9:m0_write -> mm_interconnect_0:mm_bridge_9_m0_write
	wire          mm_bridge_9_m0_read;                                           // mm_bridge_9:m0_read -> mm_interconnect_0:mm_bridge_9_m0_read
	wire  [127:0] mm_bridge_9_m0_readdata;                                       // mm_interconnect_0:mm_bridge_9_m0_readdata -> mm_bridge_9:m0_readdata
	wire          mm_bridge_9_m0_debugaccess;                                    // mm_bridge_9:m0_debugaccess -> mm_interconnect_0:mm_bridge_9_m0_debugaccess
	wire   [15:0] mm_bridge_9_m0_byteenable;                                     // mm_bridge_9:m0_byteenable -> mm_interconnect_0:mm_bridge_9_m0_byteenable
	wire          mm_bridge_9_m0_readdatavalid;                                  // mm_interconnect_0:mm_bridge_9_m0_readdatavalid -> mm_bridge_9:m0_readdatavalid
	wire    [2:0] mm_bridge_7_m0_burstcount;                                     // mm_bridge_7:m0_burstcount -> mm_interconnect_0:mm_bridge_7_m0_burstcount
	wire          mm_bridge_7_m0_waitrequest;                                    // mm_interconnect_0:mm_bridge_7_m0_waitrequest -> mm_bridge_7:m0_waitrequest
	wire   [25:0] mm_bridge_7_m0_address;                                        // mm_bridge_7:m0_address -> mm_interconnect_0:mm_bridge_7_m0_address
	wire  [127:0] mm_bridge_7_m0_writedata;                                      // mm_bridge_7:m0_writedata -> mm_interconnect_0:mm_bridge_7_m0_writedata
	wire          mm_bridge_7_m0_write;                                          // mm_bridge_7:m0_write -> mm_interconnect_0:mm_bridge_7_m0_write
	wire          mm_bridge_7_m0_read;                                           // mm_bridge_7:m0_read -> mm_interconnect_0:mm_bridge_7_m0_read
	wire  [127:0] mm_bridge_7_m0_readdata;                                       // mm_interconnect_0:mm_bridge_7_m0_readdata -> mm_bridge_7:m0_readdata
	wire          mm_bridge_7_m0_debugaccess;                                    // mm_bridge_7:m0_debugaccess -> mm_interconnect_0:mm_bridge_7_m0_debugaccess
	wire   [15:0] mm_bridge_7_m0_byteenable;                                     // mm_bridge_7:m0_byteenable -> mm_interconnect_0:mm_bridge_7_m0_byteenable
	wire          mm_bridge_7_m0_readdatavalid;                                  // mm_interconnect_0:mm_bridge_7_m0_readdatavalid -> mm_bridge_7:m0_readdatavalid
	wire    [2:0] mm_bridge_5_m0_burstcount;                                     // mm_bridge_5:m0_burstcount -> mm_interconnect_0:mm_bridge_5_m0_burstcount
	wire          mm_bridge_5_m0_waitrequest;                                    // mm_interconnect_0:mm_bridge_5_m0_waitrequest -> mm_bridge_5:m0_waitrequest
	wire   [25:0] mm_bridge_5_m0_address;                                        // mm_bridge_5:m0_address -> mm_interconnect_0:mm_bridge_5_m0_address
	wire  [127:0] mm_bridge_5_m0_writedata;                                      // mm_bridge_5:m0_writedata -> mm_interconnect_0:mm_bridge_5_m0_writedata
	wire          mm_bridge_5_m0_write;                                          // mm_bridge_5:m0_write -> mm_interconnect_0:mm_bridge_5_m0_write
	wire          mm_bridge_5_m0_read;                                           // mm_bridge_5:m0_read -> mm_interconnect_0:mm_bridge_5_m0_read
	wire  [127:0] mm_bridge_5_m0_readdata;                                       // mm_interconnect_0:mm_bridge_5_m0_readdata -> mm_bridge_5:m0_readdata
	wire          mm_bridge_5_m0_debugaccess;                                    // mm_bridge_5:m0_debugaccess -> mm_interconnect_0:mm_bridge_5_m0_debugaccess
	wire   [15:0] mm_bridge_5_m0_byteenable;                                     // mm_bridge_5:m0_byteenable -> mm_interconnect_0:mm_bridge_5_m0_byteenable
	wire          mm_bridge_5_m0_readdatavalid;                                  // mm_interconnect_0:mm_bridge_5_m0_readdatavalid -> mm_bridge_5:m0_readdatavalid
	wire    [2:0] mm_bridge_10_m0_burstcount;                                    // mm_bridge_10:m0_burstcount -> mm_interconnect_0:mm_bridge_10_m0_burstcount
	wire          mm_bridge_10_m0_waitrequest;                                   // mm_interconnect_0:mm_bridge_10_m0_waitrequest -> mm_bridge_10:m0_waitrequest
	wire   [25:0] mm_bridge_10_m0_address;                                       // mm_bridge_10:m0_address -> mm_interconnect_0:mm_bridge_10_m0_address
	wire  [127:0] mm_bridge_10_m0_writedata;                                     // mm_bridge_10:m0_writedata -> mm_interconnect_0:mm_bridge_10_m0_writedata
	wire          mm_bridge_10_m0_write;                                         // mm_bridge_10:m0_write -> mm_interconnect_0:mm_bridge_10_m0_write
	wire          mm_bridge_10_m0_read;                                          // mm_bridge_10:m0_read -> mm_interconnect_0:mm_bridge_10_m0_read
	wire  [127:0] mm_bridge_10_m0_readdata;                                      // mm_interconnect_0:mm_bridge_10_m0_readdata -> mm_bridge_10:m0_readdata
	wire          mm_bridge_10_m0_debugaccess;                                   // mm_bridge_10:m0_debugaccess -> mm_interconnect_0:mm_bridge_10_m0_debugaccess
	wire   [15:0] mm_bridge_10_m0_byteenable;                                    // mm_bridge_10:m0_byteenable -> mm_interconnect_0:mm_bridge_10_m0_byteenable
	wire          mm_bridge_10_m0_readdatavalid;                                 // mm_interconnect_0:mm_bridge_10_m0_readdatavalid -> mm_bridge_10:m0_readdatavalid
	wire    [2:0] mm_bridge_2_m0_burstcount;                                     // mm_bridge_2:m0_burstcount -> mm_interconnect_0:mm_bridge_2_m0_burstcount
	wire          mm_bridge_2_m0_waitrequest;                                    // mm_interconnect_0:mm_bridge_2_m0_waitrequest -> mm_bridge_2:m0_waitrequest
	wire   [25:0] mm_bridge_2_m0_address;                                        // mm_bridge_2:m0_address -> mm_interconnect_0:mm_bridge_2_m0_address
	wire  [127:0] mm_bridge_2_m0_writedata;                                      // mm_bridge_2:m0_writedata -> mm_interconnect_0:mm_bridge_2_m0_writedata
	wire          mm_bridge_2_m0_write;                                          // mm_bridge_2:m0_write -> mm_interconnect_0:mm_bridge_2_m0_write
	wire          mm_bridge_2_m0_read;                                           // mm_bridge_2:m0_read -> mm_interconnect_0:mm_bridge_2_m0_read
	wire  [127:0] mm_bridge_2_m0_readdata;                                       // mm_interconnect_0:mm_bridge_2_m0_readdata -> mm_bridge_2:m0_readdata
	wire          mm_bridge_2_m0_debugaccess;                                    // mm_bridge_2:m0_debugaccess -> mm_interconnect_0:mm_bridge_2_m0_debugaccess
	wire   [15:0] mm_bridge_2_m0_byteenable;                                     // mm_bridge_2:m0_byteenable -> mm_interconnect_0:mm_bridge_2_m0_byteenable
	wire          mm_bridge_2_m0_readdatavalid;                                  // mm_interconnect_0:mm_bridge_2_m0_readdatavalid -> mm_bridge_2:m0_readdatavalid
	wire    [2:0] mm_bridge_6_m0_burstcount;                                     // mm_bridge_6:m0_burstcount -> mm_interconnect_0:mm_bridge_6_m0_burstcount
	wire          mm_bridge_6_m0_waitrequest;                                    // mm_interconnect_0:mm_bridge_6_m0_waitrequest -> mm_bridge_6:m0_waitrequest
	wire   [25:0] mm_bridge_6_m0_address;                                        // mm_bridge_6:m0_address -> mm_interconnect_0:mm_bridge_6_m0_address
	wire  [127:0] mm_bridge_6_m0_writedata;                                      // mm_bridge_6:m0_writedata -> mm_interconnect_0:mm_bridge_6_m0_writedata
	wire          mm_bridge_6_m0_write;                                          // mm_bridge_6:m0_write -> mm_interconnect_0:mm_bridge_6_m0_write
	wire          mm_bridge_6_m0_read;                                           // mm_bridge_6:m0_read -> mm_interconnect_0:mm_bridge_6_m0_read
	wire  [127:0] mm_bridge_6_m0_readdata;                                       // mm_interconnect_0:mm_bridge_6_m0_readdata -> mm_bridge_6:m0_readdata
	wire          mm_bridge_6_m0_debugaccess;                                    // mm_bridge_6:m0_debugaccess -> mm_interconnect_0:mm_bridge_6_m0_debugaccess
	wire   [15:0] mm_bridge_6_m0_byteenable;                                     // mm_bridge_6:m0_byteenable -> mm_interconnect_0:mm_bridge_6_m0_byteenable
	wire          mm_bridge_6_m0_readdatavalid;                                  // mm_interconnect_0:mm_bridge_6_m0_readdatavalid -> mm_bridge_6:m0_readdatavalid
	wire    [2:0] mm_bridge_4_m0_burstcount;                                     // mm_bridge_4:m0_burstcount -> mm_interconnect_0:mm_bridge_4_m0_burstcount
	wire          mm_bridge_4_m0_waitrequest;                                    // mm_interconnect_0:mm_bridge_4_m0_waitrequest -> mm_bridge_4:m0_waitrequest
	wire   [25:0] mm_bridge_4_m0_address;                                        // mm_bridge_4:m0_address -> mm_interconnect_0:mm_bridge_4_m0_address
	wire  [127:0] mm_bridge_4_m0_writedata;                                      // mm_bridge_4:m0_writedata -> mm_interconnect_0:mm_bridge_4_m0_writedata
	wire          mm_bridge_4_m0_write;                                          // mm_bridge_4:m0_write -> mm_interconnect_0:mm_bridge_4_m0_write
	wire          mm_bridge_4_m0_read;                                           // mm_bridge_4:m0_read -> mm_interconnect_0:mm_bridge_4_m0_read
	wire  [127:0] mm_bridge_4_m0_readdata;                                       // mm_interconnect_0:mm_bridge_4_m0_readdata -> mm_bridge_4:m0_readdata
	wire          mm_bridge_4_m0_debugaccess;                                    // mm_bridge_4:m0_debugaccess -> mm_interconnect_0:mm_bridge_4_m0_debugaccess
	wire   [15:0] mm_bridge_4_m0_byteenable;                                     // mm_bridge_4:m0_byteenable -> mm_interconnect_0:mm_bridge_4_m0_byteenable
	wire          mm_bridge_4_m0_readdatavalid;                                  // mm_interconnect_0:mm_bridge_4_m0_readdatavalid -> mm_bridge_4:m0_readdatavalid
	wire    [2:0] mm_bridge_1_m0_burstcount;                                     // mm_bridge_1:m0_burstcount -> mm_interconnect_0:mm_bridge_1_m0_burstcount
	wire          mm_bridge_1_m0_waitrequest;                                    // mm_interconnect_0:mm_bridge_1_m0_waitrequest -> mm_bridge_1:m0_waitrequest
	wire   [25:0] mm_bridge_1_m0_address;                                        // mm_bridge_1:m0_address -> mm_interconnect_0:mm_bridge_1_m0_address
	wire  [127:0] mm_bridge_1_m0_writedata;                                      // mm_bridge_1:m0_writedata -> mm_interconnect_0:mm_bridge_1_m0_writedata
	wire          mm_bridge_1_m0_write;                                          // mm_bridge_1:m0_write -> mm_interconnect_0:mm_bridge_1_m0_write
	wire          mm_bridge_1_m0_read;                                           // mm_bridge_1:m0_read -> mm_interconnect_0:mm_bridge_1_m0_read
	wire  [127:0] mm_bridge_1_m0_readdata;                                       // mm_interconnect_0:mm_bridge_1_m0_readdata -> mm_bridge_1:m0_readdata
	wire          mm_bridge_1_m0_debugaccess;                                    // mm_bridge_1:m0_debugaccess -> mm_interconnect_0:mm_bridge_1_m0_debugaccess
	wire   [15:0] mm_bridge_1_m0_byteenable;                                     // mm_bridge_1:m0_byteenable -> mm_interconnect_0:mm_bridge_1_m0_byteenable
	wire          mm_bridge_1_m0_readdatavalid;                                  // mm_interconnect_0:mm_bridge_1_m0_readdatavalid -> mm_bridge_1:m0_readdatavalid
	wire    [2:0] mm_bridge_3_m0_burstcount;                                     // mm_bridge_3:m0_burstcount -> mm_interconnect_0:mm_bridge_3_m0_burstcount
	wire          mm_bridge_3_m0_waitrequest;                                    // mm_interconnect_0:mm_bridge_3_m0_waitrequest -> mm_bridge_3:m0_waitrequest
	wire   [25:0] mm_bridge_3_m0_address;                                        // mm_bridge_3:m0_address -> mm_interconnect_0:mm_bridge_3_m0_address
	wire  [127:0] mm_bridge_3_m0_writedata;                                      // mm_bridge_3:m0_writedata -> mm_interconnect_0:mm_bridge_3_m0_writedata
	wire          mm_bridge_3_m0_write;                                          // mm_bridge_3:m0_write -> mm_interconnect_0:mm_bridge_3_m0_write
	wire          mm_bridge_3_m0_read;                                           // mm_bridge_3:m0_read -> mm_interconnect_0:mm_bridge_3_m0_read
	wire  [127:0] mm_bridge_3_m0_readdata;                                       // mm_interconnect_0:mm_bridge_3_m0_readdata -> mm_bridge_3:m0_readdata
	wire          mm_bridge_3_m0_debugaccess;                                    // mm_bridge_3:m0_debugaccess -> mm_interconnect_0:mm_bridge_3_m0_debugaccess
	wire   [15:0] mm_bridge_3_m0_byteenable;                                     // mm_bridge_3:m0_byteenable -> mm_interconnect_0:mm_bridge_3_m0_byteenable
	wire          mm_bridge_3_m0_readdatavalid;                                  // mm_interconnect_0:mm_bridge_3_m0_readdatavalid -> mm_bridge_3:m0_readdatavalid
	wire    [2:0] mm_bridge_8_m0_burstcount;                                     // mm_bridge_8:m0_burstcount -> mm_interconnect_0:mm_bridge_8_m0_burstcount
	wire          mm_bridge_8_m0_waitrequest;                                    // mm_interconnect_0:mm_bridge_8_m0_waitrequest -> mm_bridge_8:m0_waitrequest
	wire   [25:0] mm_bridge_8_m0_address;                                        // mm_bridge_8:m0_address -> mm_interconnect_0:mm_bridge_8_m0_address
	wire  [127:0] mm_bridge_8_m0_writedata;                                      // mm_bridge_8:m0_writedata -> mm_interconnect_0:mm_bridge_8_m0_writedata
	wire          mm_bridge_8_m0_write;                                          // mm_bridge_8:m0_write -> mm_interconnect_0:mm_bridge_8_m0_write
	wire          mm_bridge_8_m0_read;                                           // mm_bridge_8:m0_read -> mm_interconnect_0:mm_bridge_8_m0_read
	wire  [127:0] mm_bridge_8_m0_readdata;                                       // mm_interconnect_0:mm_bridge_8_m0_readdata -> mm_bridge_8:m0_readdata
	wire          mm_bridge_8_m0_debugaccess;                                    // mm_bridge_8:m0_debugaccess -> mm_interconnect_0:mm_bridge_8_m0_debugaccess
	wire   [15:0] mm_bridge_8_m0_byteenable;                                     // mm_bridge_8:m0_byteenable -> mm_interconnect_0:mm_bridge_8_m0_byteenable
	wire          mm_bridge_8_m0_readdatavalid;                                  // mm_interconnect_0:mm_bridge_8_m0_readdatavalid -> mm_bridge_8:m0_readdatavalid
	wire    [2:0] mm_bridge_0_m0_burstcount;                                     // mm_bridge_0:m0_burstcount -> mm_interconnect_0:mm_bridge_0_m0_burstcount
	wire          mm_bridge_0_m0_waitrequest;                                    // mm_interconnect_0:mm_bridge_0_m0_waitrequest -> mm_bridge_0:m0_waitrequest
	wire   [25:0] mm_bridge_0_m0_address;                                        // mm_bridge_0:m0_address -> mm_interconnect_0:mm_bridge_0_m0_address
	wire  [127:0] mm_bridge_0_m0_writedata;                                      // mm_bridge_0:m0_writedata -> mm_interconnect_0:mm_bridge_0_m0_writedata
	wire          mm_bridge_0_m0_write;                                          // mm_bridge_0:m0_write -> mm_interconnect_0:mm_bridge_0_m0_write
	wire          mm_bridge_0_m0_read;                                           // mm_bridge_0:m0_read -> mm_interconnect_0:mm_bridge_0_m0_read
	wire  [127:0] mm_bridge_0_m0_readdata;                                       // mm_interconnect_0:mm_bridge_0_m0_readdata -> mm_bridge_0:m0_readdata
	wire          mm_bridge_0_m0_debugaccess;                                    // mm_bridge_0:m0_debugaccess -> mm_interconnect_0:mm_bridge_0_m0_debugaccess
	wire   [15:0] mm_bridge_0_m0_byteenable;                                     // mm_bridge_0:m0_byteenable -> mm_interconnect_0:mm_bridge_0_m0_byteenable
	wire          mm_bridge_0_m0_readdatavalid;                                  // mm_interconnect_0:mm_bridge_0_m0_readdatavalid -> mm_bridge_0:m0_readdatavalid
	wire          rst_controller_reset_out_reset;                                // rst_controller:reset_out -> [mm_bridge_0:reset, mm_bridge_10:reset, mm_bridge_1:reset, mm_bridge_2:reset, mm_bridge_3:reset, mm_bridge_4:reset, mm_bridge_5:reset, mm_bridge_6:reset, mm_bridge_7:reset, mm_bridge_8:reset, mm_interconnect_0:mm_bridge_0_reset_reset_bridge_in_reset_reset]
	wire          rst_controller_001_reset_out_reset;                            // rst_controller_001:reset_out -> [mm_bridge_9:reset, mm_interconnect_0:mm_bridge_9_reset_reset_bridge_in_reset_reset]
	wire          rst_controller_002_reset_out_reset;                            // rst_controller_002:reset_out -> [mm_interconnect_0:mem_if_ddr3_emif_0_avl_0_translator_reset_reset_bridge_in_reset_reset, mm_interconnect_0:mem_if_ddr3_emif_0_mp_cmd_reset_n_0_reset_bridge_in_reset_reset]

	soc_system_mem_0_mem_if_ddr3_emif_0 mem_if_ddr3_emif_0 (
		.pll_ref_clk                (clk_clk),                                                       //        pll_ref_clk.clk
		.global_reset_n             (reset_reset_n),                                                 //       global_reset.reset_n
		.soft_reset_n               (reset_reset_n),                                                 //         soft_reset.reset_n
		.afi_clk                    (mem_if_ddr3_emif_0_afi_clk_clk),                                //            afi_clk.clk
		.afi_half_clk               (afi_clk_clk),                                                   //       afi_half_clk.clk
		.afi_reset_n                (),                                                              //          afi_reset.reset_n
		.afi_reset_export_n         (),                                                              //   afi_reset_export.reset_n
		.mem_a                      (memory_0_mem_a),                                                //             memory.mem_a
		.mem_ba                     (memory_0_mem_ba),                                               //                   .mem_ba
		.mem_ck                     (memory_0_mem_ck),                                               //                   .mem_ck
		.mem_ck_n                   (memory_0_mem_ck_n),                                             //                   .mem_ck_n
		.mem_cke                    (memory_0_mem_cke),                                              //                   .mem_cke
		.mem_cs_n                   (memory_0_mem_cs_n),                                             //                   .mem_cs_n
		.mem_dm                     (memory_0_mem_dm),                                               //                   .mem_dm
		.mem_ras_n                  (memory_0_mem_ras_n),                                            //                   .mem_ras_n
		.mem_cas_n                  (memory_0_mem_cas_n),                                            //                   .mem_cas_n
		.mem_we_n                   (memory_0_mem_we_n),                                             //                   .mem_we_n
		.mem_reset_n                (memory_0_mem_reset_n),                                          //                   .mem_reset_n
		.mem_dq                     (memory_0_mem_dq),                                               //                   .mem_dq
		.mem_dqs                    (memory_0_mem_dqs),                                              //                   .mem_dqs
		.mem_dqs_n                  (memory_0_mem_dqs_n),                                            //                   .mem_dqs_n
		.mem_odt                    (memory_0_mem_odt),                                              //                   .mem_odt
		.avl_ready_0                (mm_interconnect_0_mem_if_ddr3_emif_0_avl_0_waitrequest),        //              avl_0.waitrequest_n
		.avl_burstbegin_0           (mm_interconnect_0_mem_if_ddr3_emif_0_avl_0_beginbursttransfer), //                   .beginbursttransfer
		.avl_addr_0                 (mm_interconnect_0_mem_if_ddr3_emif_0_avl_0_address),            //                   .address
		.avl_rdata_valid_0          (mm_interconnect_0_mem_if_ddr3_emif_0_avl_0_readdatavalid),      //                   .readdatavalid
		.avl_rdata_0                (mm_interconnect_0_mem_if_ddr3_emif_0_avl_0_readdata),           //                   .readdata
		.avl_wdata_0                (mm_interconnect_0_mem_if_ddr3_emif_0_avl_0_writedata),          //                   .writedata
		.avl_be_0                   (mm_interconnect_0_mem_if_ddr3_emif_0_avl_0_byteenable),         //                   .byteenable
		.avl_read_req_0             (mm_interconnect_0_mem_if_ddr3_emif_0_avl_0_read),               //                   .read
		.avl_write_req_0            (mm_interconnect_0_mem_if_ddr3_emif_0_avl_0_write),              //                   .write
		.avl_size_0                 (mm_interconnect_0_mem_if_ddr3_emif_0_avl_0_burstcount),         //                   .burstcount
		.mp_cmd_clk_0_clk           (mem_if_ddr3_emif_0_afi_clk_clk),                                //       mp_cmd_clk_0.clk
		.mp_cmd_reset_n_0_reset_n   (reset_reset_n),                                                 //   mp_cmd_reset_n_0.reset_n
		.mp_rfifo_clk_0_clk         (mem_if_ddr3_emif_0_afi_clk_clk),                                //     mp_rfifo_clk_0.clk
		.mp_rfifo_reset_n_0_reset_n (reset_reset_n),                                                 // mp_rfifo_reset_n_0.reset_n
		.mp_wfifo_clk_0_clk         (mem_if_ddr3_emif_0_afi_clk_clk),                                //     mp_wfifo_clk_0.clk
		.mp_wfifo_reset_n_0_reset_n (reset_reset_n),                                                 // mp_wfifo_reset_n_0.reset_n
		.local_init_done            (mem_if_ddr3_emif_0_status_local_init_done),                     //             status.local_init_done
		.local_cal_success          (mem_if_ddr3_emif_0_status_local_cal_success),                   //                   .local_cal_success
		.local_cal_fail             (mem_if_ddr3_emif_0_status_local_cal_fail),                      //                   .local_cal_fail
		.oct_rzqin                  (oct_rzqin),                                                     //                oct.rzqin
		.pll_mem_clk                (mem_if_ddr3_emif_0_pll_sharing_pll_mem_clk),                    //        pll_sharing.pll_mem_clk
		.pll_write_clk              (mem_if_ddr3_emif_0_pll_sharing_pll_write_clk),                  //                   .pll_write_clk
		.pll_locked                 (mem_if_ddr3_emif_0_pll_sharing_pll_locked),                     //                   .pll_locked
		.pll_write_clk_pre_phy_clk  (mem_if_ddr3_emif_0_pll_sharing_pll_write_clk_pre_phy_clk),      //                   .pll_write_clk_pre_phy_clk
		.pll_addr_cmd_clk           (mem_if_ddr3_emif_0_pll_sharing_pll_addr_cmd_clk),               //                   .pll_addr_cmd_clk
		.pll_avl_clk                (mem_if_ddr3_emif_0_pll_sharing_pll_avl_clk),                    //                   .pll_avl_clk
		.pll_config_clk             (mem_if_ddr3_emif_0_pll_sharing_pll_config_clk),                 //                   .pll_config_clk
		.pll_dr_clk                 (mem_if_ddr3_emif_0_pll_sharing_pll_dr_clk),                     //                   .pll_dr_clk
		.pll_dr_clk_pre_phy_clk     (mem_if_ddr3_emif_0_pll_sharing_pll_dr_clk_pre_phy_clk),         //                   .pll_dr_clk_pre_phy_clk
		.pll_mem_phy_clk            (mem_if_ddr3_emif_0_pll_sharing_pll_mem_phy_clk),                //                   .pll_mem_phy_clk
		.afi_phy_clk                (mem_if_ddr3_emif_0_pll_sharing_afi_phy_clk),                    //                   .afi_phy_clk
		.pll_avl_phy_clk            (mem_if_ddr3_emif_0_pll_sharing_pll_avl_phy_clk)                 //                   .pll_avl_phy_clk
	);

	altera_avalon_mm_bridge #(
		.DATA_WIDTH        (128),
		.SYMBOL_WIDTH      (8),
		.ADDRESS_WIDTH     (26),
		.BURSTCOUNT_WIDTH  (3),
		.PIPELINE_COMMAND  (1),
		.PIPELINE_RESPONSE (1)
	) mm_bridge_0 (
		.clk              (afi_clk_clk),                    //   clk.clk
		.reset            (rst_controller_reset_out_reset), // reset.reset
		.s0_waitrequest   (mem0_waitrequest),               //    s0.waitrequest
		.s0_readdata      (mem0_readdata),                  //      .readdata
		.s0_readdatavalid (mem0_readdatavalid),             //      .readdatavalid
		.s0_burstcount    (mem0_burstcount),                //      .burstcount
		.s0_writedata     (mem0_writedata),                 //      .writedata
		.s0_address       (mem0_address),                   //      .address
		.s0_write         (mem0_write),                     //      .write
		.s0_read          (mem0_read),                      //      .read
		.s0_byteenable    (mem0_byteenable),                //      .byteenable
		.s0_debugaccess   (mem0_debugaccess),               //      .debugaccess
		.m0_waitrequest   (mm_bridge_0_m0_waitrequest),     //    m0.waitrequest
		.m0_readdata      (mm_bridge_0_m0_readdata),        //      .readdata
		.m0_readdatavalid (mm_bridge_0_m0_readdatavalid),   //      .readdatavalid
		.m0_burstcount    (mm_bridge_0_m0_burstcount),      //      .burstcount
		.m0_writedata     (mm_bridge_0_m0_writedata),       //      .writedata
		.m0_address       (mm_bridge_0_m0_address),         //      .address
		.m0_write         (mm_bridge_0_m0_write),           //      .write
		.m0_read          (mm_bridge_0_m0_read),            //      .read
		.m0_byteenable    (mm_bridge_0_m0_byteenable),      //      .byteenable
		.m0_debugaccess   (mm_bridge_0_m0_debugaccess)      //      .debugaccess
	);

	altera_avalon_mm_bridge #(
		.DATA_WIDTH        (128),
		.SYMBOL_WIDTH      (8),
		.ADDRESS_WIDTH     (26),
		.BURSTCOUNT_WIDTH  (3),
		.PIPELINE_COMMAND  (1),
		.PIPELINE_RESPONSE (1)
	) mm_bridge_1 (
		.clk              (afi_clk_clk),                    //   clk.clk
		.reset            (rst_controller_reset_out_reset), // reset.reset
		.s0_waitrequest   (mem1_waitrequest),               //    s0.waitrequest
		.s0_readdata      (mem1_readdata),                  //      .readdata
		.s0_readdatavalid (mem1_readdatavalid),             //      .readdatavalid
		.s0_burstcount    (mem1_burstcount),                //      .burstcount
		.s0_writedata     (mem1_writedata),                 //      .writedata
		.s0_address       (mem1_address),                   //      .address
		.s0_write         (mem1_write),                     //      .write
		.s0_read          (mem1_read),                      //      .read
		.s0_byteenable    (mem1_byteenable),                //      .byteenable
		.s0_debugaccess   (mem1_debugaccess),               //      .debugaccess
		.m0_waitrequest   (mm_bridge_1_m0_waitrequest),     //    m0.waitrequest
		.m0_readdata      (mm_bridge_1_m0_readdata),        //      .readdata
		.m0_readdatavalid (mm_bridge_1_m0_readdatavalid),   //      .readdatavalid
		.m0_burstcount    (mm_bridge_1_m0_burstcount),      //      .burstcount
		.m0_writedata     (mm_bridge_1_m0_writedata),       //      .writedata
		.m0_address       (mm_bridge_1_m0_address),         //      .address
		.m0_write         (mm_bridge_1_m0_write),           //      .write
		.m0_read          (mm_bridge_1_m0_read),            //      .read
		.m0_byteenable    (mm_bridge_1_m0_byteenable),      //      .byteenable
		.m0_debugaccess   (mm_bridge_1_m0_debugaccess)      //      .debugaccess
	);

	altera_avalon_mm_bridge #(
		.DATA_WIDTH        (128),
		.SYMBOL_WIDTH      (8),
		.ADDRESS_WIDTH     (26),
		.BURSTCOUNT_WIDTH  (3),
		.PIPELINE_COMMAND  (1),
		.PIPELINE_RESPONSE (1)
	) mm_bridge_2 (
		.clk              (afi_clk_clk),                    //   clk.clk
		.reset            (rst_controller_reset_out_reset), // reset.reset
		.s0_waitrequest   (mem2_waitrequest),               //    s0.waitrequest
		.s0_readdata      (mem2_readdata),                  //      .readdata
		.s0_readdatavalid (mem2_readdatavalid),             //      .readdatavalid
		.s0_burstcount    (mem2_burstcount),                //      .burstcount
		.s0_writedata     (mem2_writedata),                 //      .writedata
		.s0_address       (mem2_address),                   //      .address
		.s0_write         (mem2_write),                     //      .write
		.s0_read          (mem2_read),                      //      .read
		.s0_byteenable    (mem2_byteenable),                //      .byteenable
		.s0_debugaccess   (mem2_debugaccess),               //      .debugaccess
		.m0_waitrequest   (mm_bridge_2_m0_waitrequest),     //    m0.waitrequest
		.m0_readdata      (mm_bridge_2_m0_readdata),        //      .readdata
		.m0_readdatavalid (mm_bridge_2_m0_readdatavalid),   //      .readdatavalid
		.m0_burstcount    (mm_bridge_2_m0_burstcount),      //      .burstcount
		.m0_writedata     (mm_bridge_2_m0_writedata),       //      .writedata
		.m0_address       (mm_bridge_2_m0_address),         //      .address
		.m0_write         (mm_bridge_2_m0_write),           //      .write
		.m0_read          (mm_bridge_2_m0_read),            //      .read
		.m0_byteenable    (mm_bridge_2_m0_byteenable),      //      .byteenable
		.m0_debugaccess   (mm_bridge_2_m0_debugaccess)      //      .debugaccess
	);

	altera_avalon_mm_bridge #(
		.DATA_WIDTH        (128),
		.SYMBOL_WIDTH      (8),
		.ADDRESS_WIDTH     (26),
		.BURSTCOUNT_WIDTH  (3),
		.PIPELINE_COMMAND  (1),
		.PIPELINE_RESPONSE (1)
	) mm_bridge_3 (
		.clk              (afi_clk_clk),                    //   clk.clk
		.reset            (rst_controller_reset_out_reset), // reset.reset
		.s0_waitrequest   (mem3_waitrequest),               //    s0.waitrequest
		.s0_readdata      (mem3_readdata),                  //      .readdata
		.s0_readdatavalid (mem3_readdatavalid),             //      .readdatavalid
		.s0_burstcount    (mem3_burstcount),                //      .burstcount
		.s0_writedata     (mem3_writedata),                 //      .writedata
		.s0_address       (mem3_address),                   //      .address
		.s0_write         (mem3_write),                     //      .write
		.s0_read          (mem3_read),                      //      .read
		.s0_byteenable    (mem3_byteenable),                //      .byteenable
		.s0_debugaccess   (mem3_debugaccess),               //      .debugaccess
		.m0_waitrequest   (mm_bridge_3_m0_waitrequest),     //    m0.waitrequest
		.m0_readdata      (mm_bridge_3_m0_readdata),        //      .readdata
		.m0_readdatavalid (mm_bridge_3_m0_readdatavalid),   //      .readdatavalid
		.m0_burstcount    (mm_bridge_3_m0_burstcount),      //      .burstcount
		.m0_writedata     (mm_bridge_3_m0_writedata),       //      .writedata
		.m0_address       (mm_bridge_3_m0_address),         //      .address
		.m0_write         (mm_bridge_3_m0_write),           //      .write
		.m0_read          (mm_bridge_3_m0_read),            //      .read
		.m0_byteenable    (mm_bridge_3_m0_byteenable),      //      .byteenable
		.m0_debugaccess   (mm_bridge_3_m0_debugaccess)      //      .debugaccess
	);

	altera_avalon_mm_bridge #(
		.DATA_WIDTH        (128),
		.SYMBOL_WIDTH      (8),
		.ADDRESS_WIDTH     (26),
		.BURSTCOUNT_WIDTH  (3),
		.PIPELINE_COMMAND  (1),
		.PIPELINE_RESPONSE (1)
	) mm_bridge_4 (
		.clk              (afi_clk_clk),                    //   clk.clk
		.reset            (rst_controller_reset_out_reset), // reset.reset
		.s0_waitrequest   (mem4_waitrequest),               //    s0.waitrequest
		.s0_readdata      (mem4_readdata),                  //      .readdata
		.s0_readdatavalid (mem4_readdatavalid),             //      .readdatavalid
		.s0_burstcount    (mem4_burstcount),                //      .burstcount
		.s0_writedata     (mem4_writedata),                 //      .writedata
		.s0_address       (mem4_address),                   //      .address
		.s0_write         (mem4_write),                     //      .write
		.s0_read          (mem4_read),                      //      .read
		.s0_byteenable    (mem4_byteenable),                //      .byteenable
		.s0_debugaccess   (mem4_debugaccess),               //      .debugaccess
		.m0_waitrequest   (mm_bridge_4_m0_waitrequest),     //    m0.waitrequest
		.m0_readdata      (mm_bridge_4_m0_readdata),        //      .readdata
		.m0_readdatavalid (mm_bridge_4_m0_readdatavalid),   //      .readdatavalid
		.m0_burstcount    (mm_bridge_4_m0_burstcount),      //      .burstcount
		.m0_writedata     (mm_bridge_4_m0_writedata),       //      .writedata
		.m0_address       (mm_bridge_4_m0_address),         //      .address
		.m0_write         (mm_bridge_4_m0_write),           //      .write
		.m0_read          (mm_bridge_4_m0_read),            //      .read
		.m0_byteenable    (mm_bridge_4_m0_byteenable),      //      .byteenable
		.m0_debugaccess   (mm_bridge_4_m0_debugaccess)      //      .debugaccess
	);

	altera_avalon_mm_bridge #(
		.DATA_WIDTH        (128),
		.SYMBOL_WIDTH      (8),
		.ADDRESS_WIDTH     (26),
		.BURSTCOUNT_WIDTH  (3),
		.PIPELINE_COMMAND  (1),
		.PIPELINE_RESPONSE (1)
	) mm_bridge_5 (
		.clk              (afi_clk_clk),                    //   clk.clk
		.reset            (rst_controller_reset_out_reset), // reset.reset
		.s0_waitrequest   (cam0_waitrequest),               //    s0.waitrequest
		.s0_readdata      (cam0_readdata),                  //      .readdata
		.s0_readdatavalid (cam0_readdatavalid),             //      .readdatavalid
		.s0_burstcount    (cam0_burstcount),                //      .burstcount
		.s0_writedata     (cam0_writedata),                 //      .writedata
		.s0_address       (cam0_address),                   //      .address
		.s0_write         (cam0_write),                     //      .write
		.s0_read          (cam0_read),                      //      .read
		.s0_byteenable    (cam0_byteenable),                //      .byteenable
		.s0_debugaccess   (cam0_debugaccess),               //      .debugaccess
		.m0_waitrequest   (mm_bridge_5_m0_waitrequest),     //    m0.waitrequest
		.m0_readdata      (mm_bridge_5_m0_readdata),        //      .readdata
		.m0_readdatavalid (mm_bridge_5_m0_readdatavalid),   //      .readdatavalid
		.m0_burstcount    (mm_bridge_5_m0_burstcount),      //      .burstcount
		.m0_writedata     (mm_bridge_5_m0_writedata),       //      .writedata
		.m0_address       (mm_bridge_5_m0_address),         //      .address
		.m0_write         (mm_bridge_5_m0_write),           //      .write
		.m0_read          (mm_bridge_5_m0_read),            //      .read
		.m0_byteenable    (mm_bridge_5_m0_byteenable),      //      .byteenable
		.m0_debugaccess   (mm_bridge_5_m0_debugaccess)      //      .debugaccess
	);

	altera_avalon_mm_bridge #(
		.DATA_WIDTH        (128),
		.SYMBOL_WIDTH      (8),
		.ADDRESS_WIDTH     (26),
		.BURSTCOUNT_WIDTH  (3),
		.PIPELINE_COMMAND  (1),
		.PIPELINE_RESPONSE (1)
	) mm_bridge_6 (
		.clk              (afi_clk_clk),                    //   clk.clk
		.reset            (rst_controller_reset_out_reset), // reset.reset
		.s0_waitrequest   (cam1_waitrequest),               //    s0.waitrequest
		.s0_readdata      (cam1_readdata),                  //      .readdata
		.s0_readdatavalid (cam1_readdatavalid),             //      .readdatavalid
		.s0_burstcount    (cam1_burstcount),                //      .burstcount
		.s0_writedata     (cam1_writedata),                 //      .writedata
		.s0_address       (cam1_address),                   //      .address
		.s0_write         (cam1_write),                     //      .write
		.s0_read          (cam1_read),                      //      .read
		.s0_byteenable    (cam1_byteenable),                //      .byteenable
		.s0_debugaccess   (cam1_debugaccess),               //      .debugaccess
		.m0_waitrequest   (mm_bridge_6_m0_waitrequest),     //    m0.waitrequest
		.m0_readdata      (mm_bridge_6_m0_readdata),        //      .readdata
		.m0_readdatavalid (mm_bridge_6_m0_readdatavalid),   //      .readdatavalid
		.m0_burstcount    (mm_bridge_6_m0_burstcount),      //      .burstcount
		.m0_writedata     (mm_bridge_6_m0_writedata),       //      .writedata
		.m0_address       (mm_bridge_6_m0_address),         //      .address
		.m0_write         (mm_bridge_6_m0_write),           //      .write
		.m0_read          (mm_bridge_6_m0_read),            //      .read
		.m0_byteenable    (mm_bridge_6_m0_byteenable),      //      .byteenable
		.m0_debugaccess   (mm_bridge_6_m0_debugaccess)      //      .debugaccess
	);

	altera_avalon_mm_bridge #(
		.DATA_WIDTH        (128),
		.SYMBOL_WIDTH      (8),
		.ADDRESS_WIDTH     (26),
		.BURSTCOUNT_WIDTH  (3),
		.PIPELINE_COMMAND  (1),
		.PIPELINE_RESPONSE (1)
	) mm_bridge_7 (
		.clk              (afi_clk_clk),                    //   clk.clk
		.reset            (rst_controller_reset_out_reset), // reset.reset
		.s0_waitrequest   (cam23_waitrequest),              //    s0.waitrequest
		.s0_readdata      (cam23_readdata),                 //      .readdata
		.s0_readdatavalid (cam23_readdatavalid),            //      .readdatavalid
		.s0_burstcount    (cam23_burstcount),               //      .burstcount
		.s0_writedata     (cam23_writedata),                //      .writedata
		.s0_address       (cam23_address),                  //      .address
		.s0_write         (cam23_write),                    //      .write
		.s0_read          (cam23_read),                     //      .read
		.s0_byteenable    (cam23_byteenable),               //      .byteenable
		.s0_debugaccess   (cam23_debugaccess),              //      .debugaccess
		.m0_waitrequest   (mm_bridge_7_m0_waitrequest),     //    m0.waitrequest
		.m0_readdata      (mm_bridge_7_m0_readdata),        //      .readdata
		.m0_readdatavalid (mm_bridge_7_m0_readdatavalid),   //      .readdatavalid
		.m0_burstcount    (mm_bridge_7_m0_burstcount),      //      .burstcount
		.m0_writedata     (mm_bridge_7_m0_writedata),       //      .writedata
		.m0_address       (mm_bridge_7_m0_address),         //      .address
		.m0_write         (mm_bridge_7_m0_write),           //      .write
		.m0_read          (mm_bridge_7_m0_read),            //      .read
		.m0_byteenable    (mm_bridge_7_m0_byteenable),      //      .byteenable
		.m0_debugaccess   (mm_bridge_7_m0_debugaccess)      //      .debugaccess
	);

	altera_avalon_mm_bridge #(
		.DATA_WIDTH        (128),
		.SYMBOL_WIDTH      (8),
		.ADDRESS_WIDTH     (26),
		.BURSTCOUNT_WIDTH  (3),
		.PIPELINE_COMMAND  (1),
		.PIPELINE_RESPONSE (1)
	) mm_bridge_8 (
		.clk              (afi_clk_clk),                    //   clk.clk
		.reset            (rst_controller_reset_out_reset), // reset.reset
		.s0_waitrequest   (cam45_waitrequest),              //    s0.waitrequest
		.s0_readdata      (cam45_readdata),                 //      .readdata
		.s0_readdatavalid (cam45_readdatavalid),            //      .readdatavalid
		.s0_burstcount    (cam45_burstcount),               //      .burstcount
		.s0_writedata     (cam45_writedata),                //      .writedata
		.s0_address       (cam45_address),                  //      .address
		.s0_write         (cam45_write),                    //      .write
		.s0_read          (cam45_read),                     //      .read
		.s0_byteenable    (cam45_byteenable),               //      .byteenable
		.s0_debugaccess   (cam45_debugaccess),              //      .debugaccess
		.m0_waitrequest   (mm_bridge_8_m0_waitrequest),     //    m0.waitrequest
		.m0_readdata      (mm_bridge_8_m0_readdata),        //      .readdata
		.m0_readdatavalid (mm_bridge_8_m0_readdatavalid),   //      .readdatavalid
		.m0_burstcount    (mm_bridge_8_m0_burstcount),      //      .burstcount
		.m0_writedata     (mm_bridge_8_m0_writedata),       //      .writedata
		.m0_address       (mm_bridge_8_m0_address),         //      .address
		.m0_write         (mm_bridge_8_m0_write),           //      .write
		.m0_read          (mm_bridge_8_m0_read),            //      .read
		.m0_byteenable    (mm_bridge_8_m0_byteenable),      //      .byteenable
		.m0_debugaccess   (mm_bridge_8_m0_debugaccess)      //      .debugaccess
	);

	altera_avalon_mm_bridge #(
		.DATA_WIDTH        (128),
		.SYMBOL_WIDTH      (8),
		.ADDRESS_WIDTH     (26),
		.BURSTCOUNT_WIDTH  (3),
		.PIPELINE_COMMAND  (1),
		.PIPELINE_RESPONSE (1)
	) mm_bridge_9 (
		.clk              (clk_0_clk),                          //   clk.clk
		.reset            (rst_controller_001_reset_out_reset), // reset.reset
		.s0_waitrequest   (hps_waitrequest),                    //    s0.waitrequest
		.s0_readdata      (hps_readdata),                       //      .readdata
		.s0_readdatavalid (hps_readdatavalid),                  //      .readdatavalid
		.s0_burstcount    (hps_burstcount),                     //      .burstcount
		.s0_writedata     (hps_writedata),                      //      .writedata
		.s0_address       (hps_address),                        //      .address
		.s0_write         (hps_write),                          //      .write
		.s0_read          (hps_read),                           //      .read
		.s0_byteenable    (hps_byteenable),                     //      .byteenable
		.s0_debugaccess   (hps_debugaccess),                    //      .debugaccess
		.m0_waitrequest   (mm_bridge_9_m0_waitrequest),         //    m0.waitrequest
		.m0_readdata      (mm_bridge_9_m0_readdata),            //      .readdata
		.m0_readdatavalid (mm_bridge_9_m0_readdatavalid),       //      .readdatavalid
		.m0_burstcount    (mm_bridge_9_m0_burstcount),          //      .burstcount
		.m0_writedata     (mm_bridge_9_m0_writedata),           //      .writedata
		.m0_address       (mm_bridge_9_m0_address),             //      .address
		.m0_write         (mm_bridge_9_m0_write),               //      .write
		.m0_read          (mm_bridge_9_m0_read),                //      .read
		.m0_byteenable    (mm_bridge_9_m0_byteenable),          //      .byteenable
		.m0_debugaccess   (mm_bridge_9_m0_debugaccess)          //      .debugaccess
	);

	altera_avalon_mm_bridge #(
		.DATA_WIDTH        (128),
		.SYMBOL_WIDTH      (8),
		.ADDRESS_WIDTH     (26),
		.BURSTCOUNT_WIDTH  (3),
		.PIPELINE_COMMAND  (1),
		.PIPELINE_RESPONSE (1)
	) mm_bridge_10 (
		.clk              (afi_clk_clk),                    //   clk.clk
		.reset            (rst_controller_reset_out_reset), // reset.reset
		.s0_waitrequest   (test_vga_waitrequest),           //    s0.waitrequest
		.s0_readdata      (test_vga_readdata),              //      .readdata
		.s0_readdatavalid (test_vga_readdatavalid),         //      .readdatavalid
		.s0_burstcount    (test_vga_burstcount),            //      .burstcount
		.s0_writedata     (test_vga_writedata),             //      .writedata
		.s0_address       (test_vga_address),               //      .address
		.s0_write         (test_vga_write),                 //      .write
		.s0_read          (test_vga_read),                  //      .read
		.s0_byteenable    (test_vga_byteenable),            //      .byteenable
		.s0_debugaccess   (test_vga_debugaccess),           //      .debugaccess
		.m0_waitrequest   (mm_bridge_10_m0_waitrequest),    //    m0.waitrequest
		.m0_readdata      (mm_bridge_10_m0_readdata),       //      .readdata
		.m0_readdatavalid (mm_bridge_10_m0_readdatavalid),  //      .readdatavalid
		.m0_burstcount    (mm_bridge_10_m0_burstcount),     //      .burstcount
		.m0_writedata     (mm_bridge_10_m0_writedata),      //      .writedata
		.m0_address       (mm_bridge_10_m0_address),        //      .address
		.m0_write         (mm_bridge_10_m0_write),          //      .write
		.m0_read          (mm_bridge_10_m0_read),           //      .read
		.m0_byteenable    (mm_bridge_10_m0_byteenable),     //      .byteenable
		.m0_debugaccess   (mm_bridge_10_m0_debugaccess)     //      .debugaccess
	);

	soc_system_mem_0_mm_interconnect_0 mm_interconnect_0 (
		.clk_1_clk_clk                                                         (clk_0_clk),                                                     //                                                       clk_1_clk.clk
		.mem_if_ddr3_emif_0_afi_clk_clk                                        (mem_if_ddr3_emif_0_afi_clk_clk),                                //                                      mem_if_ddr3_emif_0_afi_clk.clk
		.mem_if_ddr3_emif_0_afi_half_clk_clk                                   (afi_clk_clk),                                                   //                                 mem_if_ddr3_emif_0_afi_half_clk.clk
		.mem_if_ddr3_emif_0_avl_0_translator_reset_reset_bridge_in_reset_reset (rst_controller_002_reset_out_reset),                            // mem_if_ddr3_emif_0_avl_0_translator_reset_reset_bridge_in_reset.reset
		.mem_if_ddr3_emif_0_mp_cmd_reset_n_0_reset_bridge_in_reset_reset       (rst_controller_002_reset_out_reset),                            //       mem_if_ddr3_emif_0_mp_cmd_reset_n_0_reset_bridge_in_reset.reset
		.mm_bridge_0_reset_reset_bridge_in_reset_reset                         (rst_controller_reset_out_reset),                                //                         mm_bridge_0_reset_reset_bridge_in_reset.reset
		.mm_bridge_9_reset_reset_bridge_in_reset_reset                         (rst_controller_001_reset_out_reset),                            //                         mm_bridge_9_reset_reset_bridge_in_reset.reset
		.mm_bridge_0_m0_address                                                (mm_bridge_0_m0_address),                                        //                                                  mm_bridge_0_m0.address
		.mm_bridge_0_m0_waitrequest                                            (mm_bridge_0_m0_waitrequest),                                    //                                                                .waitrequest
		.mm_bridge_0_m0_burstcount                                             (mm_bridge_0_m0_burstcount),                                     //                                                                .burstcount
		.mm_bridge_0_m0_byteenable                                             (mm_bridge_0_m0_byteenable),                                     //                                                                .byteenable
		.mm_bridge_0_m0_read                                                   (mm_bridge_0_m0_read),                                           //                                                                .read
		.mm_bridge_0_m0_readdata                                               (mm_bridge_0_m0_readdata),                                       //                                                                .readdata
		.mm_bridge_0_m0_readdatavalid                                          (mm_bridge_0_m0_readdatavalid),                                  //                                                                .readdatavalid
		.mm_bridge_0_m0_write                                                  (mm_bridge_0_m0_write),                                          //                                                                .write
		.mm_bridge_0_m0_writedata                                              (mm_bridge_0_m0_writedata),                                      //                                                                .writedata
		.mm_bridge_0_m0_debugaccess                                            (mm_bridge_0_m0_debugaccess),                                    //                                                                .debugaccess
		.mm_bridge_1_m0_address                                                (mm_bridge_1_m0_address),                                        //                                                  mm_bridge_1_m0.address
		.mm_bridge_1_m0_waitrequest                                            (mm_bridge_1_m0_waitrequest),                                    //                                                                .waitrequest
		.mm_bridge_1_m0_burstcount                                             (mm_bridge_1_m0_burstcount),                                     //                                                                .burstcount
		.mm_bridge_1_m0_byteenable                                             (mm_bridge_1_m0_byteenable),                                     //                                                                .byteenable
		.mm_bridge_1_m0_read                                                   (mm_bridge_1_m0_read),                                           //                                                                .read
		.mm_bridge_1_m0_readdata                                               (mm_bridge_1_m0_readdata),                                       //                                                                .readdata
		.mm_bridge_1_m0_readdatavalid                                          (mm_bridge_1_m0_readdatavalid),                                  //                                                                .readdatavalid
		.mm_bridge_1_m0_write                                                  (mm_bridge_1_m0_write),                                          //                                                                .write
		.mm_bridge_1_m0_writedata                                              (mm_bridge_1_m0_writedata),                                      //                                                                .writedata
		.mm_bridge_1_m0_debugaccess                                            (mm_bridge_1_m0_debugaccess),                                    //                                                                .debugaccess
		.mm_bridge_10_m0_address                                               (mm_bridge_10_m0_address),                                       //                                                 mm_bridge_10_m0.address
		.mm_bridge_10_m0_waitrequest                                           (mm_bridge_10_m0_waitrequest),                                   //                                                                .waitrequest
		.mm_bridge_10_m0_burstcount                                            (mm_bridge_10_m0_burstcount),                                    //                                                                .burstcount
		.mm_bridge_10_m0_byteenable                                            (mm_bridge_10_m0_byteenable),                                    //                                                                .byteenable
		.mm_bridge_10_m0_read                                                  (mm_bridge_10_m0_read),                                          //                                                                .read
		.mm_bridge_10_m0_readdata                                              (mm_bridge_10_m0_readdata),                                      //                                                                .readdata
		.mm_bridge_10_m0_readdatavalid                                         (mm_bridge_10_m0_readdatavalid),                                 //                                                                .readdatavalid
		.mm_bridge_10_m0_write                                                 (mm_bridge_10_m0_write),                                         //                                                                .write
		.mm_bridge_10_m0_writedata                                             (mm_bridge_10_m0_writedata),                                     //                                                                .writedata
		.mm_bridge_10_m0_debugaccess                                           (mm_bridge_10_m0_debugaccess),                                   //                                                                .debugaccess
		.mm_bridge_2_m0_address                                                (mm_bridge_2_m0_address),                                        //                                                  mm_bridge_2_m0.address
		.mm_bridge_2_m0_waitrequest                                            (mm_bridge_2_m0_waitrequest),                                    //                                                                .waitrequest
		.mm_bridge_2_m0_burstcount                                             (mm_bridge_2_m0_burstcount),                                     //                                                                .burstcount
		.mm_bridge_2_m0_byteenable                                             (mm_bridge_2_m0_byteenable),                                     //                                                                .byteenable
		.mm_bridge_2_m0_read                                                   (mm_bridge_2_m0_read),                                           //                                                                .read
		.mm_bridge_2_m0_readdata                                               (mm_bridge_2_m0_readdata),                                       //                                                                .readdata
		.mm_bridge_2_m0_readdatavalid                                          (mm_bridge_2_m0_readdatavalid),                                  //                                                                .readdatavalid
		.mm_bridge_2_m0_write                                                  (mm_bridge_2_m0_write),                                          //                                                                .write
		.mm_bridge_2_m0_writedata                                              (mm_bridge_2_m0_writedata),                                      //                                                                .writedata
		.mm_bridge_2_m0_debugaccess                                            (mm_bridge_2_m0_debugaccess),                                    //                                                                .debugaccess
		.mm_bridge_3_m0_address                                                (mm_bridge_3_m0_address),                                        //                                                  mm_bridge_3_m0.address
		.mm_bridge_3_m0_waitrequest                                            (mm_bridge_3_m0_waitrequest),                                    //                                                                .waitrequest
		.mm_bridge_3_m0_burstcount                                             (mm_bridge_3_m0_burstcount),                                     //                                                                .burstcount
		.mm_bridge_3_m0_byteenable                                             (mm_bridge_3_m0_byteenable),                                     //                                                                .byteenable
		.mm_bridge_3_m0_read                                                   (mm_bridge_3_m0_read),                                           //                                                                .read
		.mm_bridge_3_m0_readdata                                               (mm_bridge_3_m0_readdata),                                       //                                                                .readdata
		.mm_bridge_3_m0_readdatavalid                                          (mm_bridge_3_m0_readdatavalid),                                  //                                                                .readdatavalid
		.mm_bridge_3_m0_write                                                  (mm_bridge_3_m0_write),                                          //                                                                .write
		.mm_bridge_3_m0_writedata                                              (mm_bridge_3_m0_writedata),                                      //                                                                .writedata
		.mm_bridge_3_m0_debugaccess                                            (mm_bridge_3_m0_debugaccess),                                    //                                                                .debugaccess
		.mm_bridge_4_m0_address                                                (mm_bridge_4_m0_address),                                        //                                                  mm_bridge_4_m0.address
		.mm_bridge_4_m0_waitrequest                                            (mm_bridge_4_m0_waitrequest),                                    //                                                                .waitrequest
		.mm_bridge_4_m0_burstcount                                             (mm_bridge_4_m0_burstcount),                                     //                                                                .burstcount
		.mm_bridge_4_m0_byteenable                                             (mm_bridge_4_m0_byteenable),                                     //                                                                .byteenable
		.mm_bridge_4_m0_read                                                   (mm_bridge_4_m0_read),                                           //                                                                .read
		.mm_bridge_4_m0_readdata                                               (mm_bridge_4_m0_readdata),                                       //                                                                .readdata
		.mm_bridge_4_m0_readdatavalid                                          (mm_bridge_4_m0_readdatavalid),                                  //                                                                .readdatavalid
		.mm_bridge_4_m0_write                                                  (mm_bridge_4_m0_write),                                          //                                                                .write
		.mm_bridge_4_m0_writedata                                              (mm_bridge_4_m0_writedata),                                      //                                                                .writedata
		.mm_bridge_4_m0_debugaccess                                            (mm_bridge_4_m0_debugaccess),                                    //                                                                .debugaccess
		.mm_bridge_5_m0_address                                                (mm_bridge_5_m0_address),                                        //                                                  mm_bridge_5_m0.address
		.mm_bridge_5_m0_waitrequest                                            (mm_bridge_5_m0_waitrequest),                                    //                                                                .waitrequest
		.mm_bridge_5_m0_burstcount                                             (mm_bridge_5_m0_burstcount),                                     //                                                                .burstcount
		.mm_bridge_5_m0_byteenable                                             (mm_bridge_5_m0_byteenable),                                     //                                                                .byteenable
		.mm_bridge_5_m0_read                                                   (mm_bridge_5_m0_read),                                           //                                                                .read
		.mm_bridge_5_m0_readdata                                               (mm_bridge_5_m0_readdata),                                       //                                                                .readdata
		.mm_bridge_5_m0_readdatavalid                                          (mm_bridge_5_m0_readdatavalid),                                  //                                                                .readdatavalid
		.mm_bridge_5_m0_write                                                  (mm_bridge_5_m0_write),                                          //                                                                .write
		.mm_bridge_5_m0_writedata                                              (mm_bridge_5_m0_writedata),                                      //                                                                .writedata
		.mm_bridge_5_m0_debugaccess                                            (mm_bridge_5_m0_debugaccess),                                    //                                                                .debugaccess
		.mm_bridge_6_m0_address                                                (mm_bridge_6_m0_address),                                        //                                                  mm_bridge_6_m0.address
		.mm_bridge_6_m0_waitrequest                                            (mm_bridge_6_m0_waitrequest),                                    //                                                                .waitrequest
		.mm_bridge_6_m0_burstcount                                             (mm_bridge_6_m0_burstcount),                                     //                                                                .burstcount
		.mm_bridge_6_m0_byteenable                                             (mm_bridge_6_m0_byteenable),                                     //                                                                .byteenable
		.mm_bridge_6_m0_read                                                   (mm_bridge_6_m0_read),                                           //                                                                .read
		.mm_bridge_6_m0_readdata                                               (mm_bridge_6_m0_readdata),                                       //                                                                .readdata
		.mm_bridge_6_m0_readdatavalid                                          (mm_bridge_6_m0_readdatavalid),                                  //                                                                .readdatavalid
		.mm_bridge_6_m0_write                                                  (mm_bridge_6_m0_write),                                          //                                                                .write
		.mm_bridge_6_m0_writedata                                              (mm_bridge_6_m0_writedata),                                      //                                                                .writedata
		.mm_bridge_6_m0_debugaccess                                            (mm_bridge_6_m0_debugaccess),                                    //                                                                .debugaccess
		.mm_bridge_7_m0_address                                                (mm_bridge_7_m0_address),                                        //                                                  mm_bridge_7_m0.address
		.mm_bridge_7_m0_waitrequest                                            (mm_bridge_7_m0_waitrequest),                                    //                                                                .waitrequest
		.mm_bridge_7_m0_burstcount                                             (mm_bridge_7_m0_burstcount),                                     //                                                                .burstcount
		.mm_bridge_7_m0_byteenable                                             (mm_bridge_7_m0_byteenable),                                     //                                                                .byteenable
		.mm_bridge_7_m0_read                                                   (mm_bridge_7_m0_read),                                           //                                                                .read
		.mm_bridge_7_m0_readdata                                               (mm_bridge_7_m0_readdata),                                       //                                                                .readdata
		.mm_bridge_7_m0_readdatavalid                                          (mm_bridge_7_m0_readdatavalid),                                  //                                                                .readdatavalid
		.mm_bridge_7_m0_write                                                  (mm_bridge_7_m0_write),                                          //                                                                .write
		.mm_bridge_7_m0_writedata                                              (mm_bridge_7_m0_writedata),                                      //                                                                .writedata
		.mm_bridge_7_m0_debugaccess                                            (mm_bridge_7_m0_debugaccess),                                    //                                                                .debugaccess
		.mm_bridge_8_m0_address                                                (mm_bridge_8_m0_address),                                        //                                                  mm_bridge_8_m0.address
		.mm_bridge_8_m0_waitrequest                                            (mm_bridge_8_m0_waitrequest),                                    //                                                                .waitrequest
		.mm_bridge_8_m0_burstcount                                             (mm_bridge_8_m0_burstcount),                                     //                                                                .burstcount
		.mm_bridge_8_m0_byteenable                                             (mm_bridge_8_m0_byteenable),                                     //                                                                .byteenable
		.mm_bridge_8_m0_read                                                   (mm_bridge_8_m0_read),                                           //                                                                .read
		.mm_bridge_8_m0_readdata                                               (mm_bridge_8_m0_readdata),                                       //                                                                .readdata
		.mm_bridge_8_m0_readdatavalid                                          (mm_bridge_8_m0_readdatavalid),                                  //                                                                .readdatavalid
		.mm_bridge_8_m0_write                                                  (mm_bridge_8_m0_write),                                          //                                                                .write
		.mm_bridge_8_m0_writedata                                              (mm_bridge_8_m0_writedata),                                      //                                                                .writedata
		.mm_bridge_8_m0_debugaccess                                            (mm_bridge_8_m0_debugaccess),                                    //                                                                .debugaccess
		.mm_bridge_9_m0_address                                                (mm_bridge_9_m0_address),                                        //                                                  mm_bridge_9_m0.address
		.mm_bridge_9_m0_waitrequest                                            (mm_bridge_9_m0_waitrequest),                                    //                                                                .waitrequest
		.mm_bridge_9_m0_burstcount                                             (mm_bridge_9_m0_burstcount),                                     //                                                                .burstcount
		.mm_bridge_9_m0_byteenable                                             (mm_bridge_9_m0_byteenable),                                     //                                                                .byteenable
		.mm_bridge_9_m0_read                                                   (mm_bridge_9_m0_read),                                           //                                                                .read
		.mm_bridge_9_m0_readdata                                               (mm_bridge_9_m0_readdata),                                       //                                                                .readdata
		.mm_bridge_9_m0_readdatavalid                                          (mm_bridge_9_m0_readdatavalid),                                  //                                                                .readdatavalid
		.mm_bridge_9_m0_write                                                  (mm_bridge_9_m0_write),                                          //                                                                .write
		.mm_bridge_9_m0_writedata                                              (mm_bridge_9_m0_writedata),                                      //                                                                .writedata
		.mm_bridge_9_m0_debugaccess                                            (mm_bridge_9_m0_debugaccess),                                    //                                                                .debugaccess
		.mem_if_ddr3_emif_0_avl_0_address                                      (mm_interconnect_0_mem_if_ddr3_emif_0_avl_0_address),            //                                        mem_if_ddr3_emif_0_avl_0.address
		.mem_if_ddr3_emif_0_avl_0_write                                        (mm_interconnect_0_mem_if_ddr3_emif_0_avl_0_write),              //                                                                .write
		.mem_if_ddr3_emif_0_avl_0_read                                         (mm_interconnect_0_mem_if_ddr3_emif_0_avl_0_read),               //                                                                .read
		.mem_if_ddr3_emif_0_avl_0_readdata                                     (mm_interconnect_0_mem_if_ddr3_emif_0_avl_0_readdata),           //                                                                .readdata
		.mem_if_ddr3_emif_0_avl_0_writedata                                    (mm_interconnect_0_mem_if_ddr3_emif_0_avl_0_writedata),          //                                                                .writedata
		.mem_if_ddr3_emif_0_avl_0_beginbursttransfer                           (mm_interconnect_0_mem_if_ddr3_emif_0_avl_0_beginbursttransfer), //                                                                .beginbursttransfer
		.mem_if_ddr3_emif_0_avl_0_burstcount                                   (mm_interconnect_0_mem_if_ddr3_emif_0_avl_0_burstcount),         //                                                                .burstcount
		.mem_if_ddr3_emif_0_avl_0_byteenable                                   (mm_interconnect_0_mem_if_ddr3_emif_0_avl_0_byteenable),         //                                                                .byteenable
		.mem_if_ddr3_emif_0_avl_0_readdatavalid                                (mm_interconnect_0_mem_if_ddr3_emif_0_avl_0_readdatavalid),      //                                                                .readdatavalid
		.mem_if_ddr3_emif_0_avl_0_waitrequest                                  (~mm_interconnect_0_mem_if_ddr3_emif_0_avl_0_waitrequest)        //                                                                .waitrequest
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                 // reset_in0.reset
		.clk            (afi_clk_clk),                    //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (clk_0_clk),                          //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (mem_if_ddr3_emif_0_afi_clk_clk),     //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
