// fpga_mem_tb.v

// Generated using ACDS version 13.1 162 at 2015.06.22.09:15:33

`timescale 1 ps / 1 ps
module fpga_mem_tb (
	);

	wire          fpga_mem_inst_clk_bfm_clk_clk;                                          // fpga_mem_inst_clk_bfm:clk -> [fpga_mem_inst:clk_clk, fpga_mem_inst_reset_bfm:clk]
	wire          fpga_mem_inst_reset_bfm_reset_reset;                                    // fpga_mem_inst_reset_bfm:reset -> [fpga_mem_inst:reset_reset_n, rst_controller:reset_in0]
	wire    [0:0] fpga_mem_inst_oct_bfm_conduit_rzqin;                                    // fpga_mem_inst_oct_bfm:sig_rzqin -> fpga_mem_inst:oct_rzqin
	wire          fpga_mem_inst_mem_if_ddr3_emif_0_status_local_cal_fail;                 // fpga_mem_inst:mem_if_ddr3_emif_0_status_local_cal_fail -> fpga_mem_inst_mem_if_ddr3_emif_0_status_bfm:sig_local_cal_fail
	wire          fpga_mem_inst_mem_if_ddr3_emif_0_status_local_cal_success;              // fpga_mem_inst:mem_if_ddr3_emif_0_status_local_cal_success -> fpga_mem_inst_mem_if_ddr3_emif_0_status_bfm:sig_local_cal_success
	wire          fpga_mem_inst_mem_if_ddr3_emif_0_status_local_init_done;                // fpga_mem_inst:mem_if_ddr3_emif_0_status_local_init_done -> fpga_mem_inst_mem_if_ddr3_emif_0_status_bfm:sig_local_init_done
	wire          fpga_mem_inst_mem_if_ddr3_emif_0_pll_sharing_pll_mem_phy_clk;           // fpga_mem_inst:mem_if_ddr3_emif_0_pll_sharing_pll_mem_phy_clk -> fpga_mem_inst_mem_if_ddr3_emif_0_pll_sharing_bfm:sig_pll_mem_phy_clk
	wire          fpga_mem_inst_mem_if_ddr3_emif_0_pll_sharing_pll_dr_clk_pre_phy_clk;    // fpga_mem_inst:mem_if_ddr3_emif_0_pll_sharing_pll_dr_clk_pre_phy_clk -> fpga_mem_inst_mem_if_ddr3_emif_0_pll_sharing_bfm:sig_pll_dr_clk_pre_phy_clk
	wire          fpga_mem_inst_mem_if_ddr3_emif_0_pll_sharing_pll_avl_clk;               // fpga_mem_inst:mem_if_ddr3_emif_0_pll_sharing_pll_avl_clk -> fpga_mem_inst_mem_if_ddr3_emif_0_pll_sharing_bfm:sig_pll_avl_clk
	wire          fpga_mem_inst_mem_if_ddr3_emif_0_pll_sharing_pll_avl_phy_clk;           // fpga_mem_inst:mem_if_ddr3_emif_0_pll_sharing_pll_avl_phy_clk -> fpga_mem_inst_mem_if_ddr3_emif_0_pll_sharing_bfm:sig_pll_avl_phy_clk
	wire          fpga_mem_inst_mem_if_ddr3_emif_0_pll_sharing_afi_phy_clk;               // fpga_mem_inst:mem_if_ddr3_emif_0_pll_sharing_afi_phy_clk -> fpga_mem_inst_mem_if_ddr3_emif_0_pll_sharing_bfm:sig_afi_phy_clk
	wire          fpga_mem_inst_mem_if_ddr3_emif_0_pll_sharing_pll_config_clk;            // fpga_mem_inst:mem_if_ddr3_emif_0_pll_sharing_pll_config_clk -> fpga_mem_inst_mem_if_ddr3_emif_0_pll_sharing_bfm:sig_pll_config_clk
	wire          fpga_mem_inst_mem_if_ddr3_emif_0_pll_sharing_pll_addr_cmd_clk;          // fpga_mem_inst:mem_if_ddr3_emif_0_pll_sharing_pll_addr_cmd_clk -> fpga_mem_inst_mem_if_ddr3_emif_0_pll_sharing_bfm:sig_pll_addr_cmd_clk
	wire          fpga_mem_inst_mem_if_ddr3_emif_0_pll_sharing_pll_dr_clk;                // fpga_mem_inst:mem_if_ddr3_emif_0_pll_sharing_pll_dr_clk -> fpga_mem_inst_mem_if_ddr3_emif_0_pll_sharing_bfm:sig_pll_dr_clk
	wire          fpga_mem_inst_mem_if_ddr3_emif_0_pll_sharing_pll_mem_clk;               // fpga_mem_inst:mem_if_ddr3_emif_0_pll_sharing_pll_mem_clk -> fpga_mem_inst_mem_if_ddr3_emif_0_pll_sharing_bfm:sig_pll_mem_clk
	wire          fpga_mem_inst_mem_if_ddr3_emif_0_pll_sharing_pll_locked;                // fpga_mem_inst:mem_if_ddr3_emif_0_pll_sharing_pll_locked -> fpga_mem_inst_mem_if_ddr3_emif_0_pll_sharing_bfm:sig_pll_locked
	wire          fpga_mem_inst_mem_if_ddr3_emif_0_pll_sharing_pll_write_clk_pre_phy_clk; // fpga_mem_inst:mem_if_ddr3_emif_0_pll_sharing_pll_write_clk_pre_phy_clk -> fpga_mem_inst_mem_if_ddr3_emif_0_pll_sharing_bfm:sig_pll_write_clk_pre_phy_clk
	wire          fpga_mem_inst_mem_if_ddr3_emif_0_pll_sharing_pll_write_clk;             // fpga_mem_inst:mem_if_ddr3_emif_0_pll_sharing_pll_write_clk -> fpga_mem_inst_mem_if_ddr3_emif_0_pll_sharing_bfm:sig_pll_write_clk
	wire          fpga_mem_inst_afi_clk_clk;                                              // fpga_mem_inst:afi_clk_clk -> [fpga_mem_inst_hps_bfm:clk, fpga_mem_inst_mr0_bfm:clk, fpga_mem_inst_mr1_bfm:clk, fpga_mem_inst_mr2_bfm:clk, fpga_mem_inst_mr3_bfm:clk, fpga_mem_inst_mrx_bfm:clk, fpga_mem_inst_mw0_bfm:clk, fpga_mem_inst_mw1_bfm:clk, fpga_mem_inst_mw2_bfm:clk, fpga_mem_inst_mw3_bfm:clk, fpga_mem_inst_mwx_bfm:clk, rst_controller:clk]
	wire          fpga_mem_inst_mrx_bfm_m0_waitrequest;                                   // fpga_mem_inst:mrx_waitrequest -> fpga_mem_inst_mrx_bfm:avm_waitrequest
	wire    [5:0] fpga_mem_inst_mrx_bfm_m0_burstcount;                                    // fpga_mem_inst_mrx_bfm:avm_burstcount -> fpga_mem_inst:mrx_burstcount
	wire  [127:0] fpga_mem_inst_mrx_bfm_m0_writedata;                                     // fpga_mem_inst_mrx_bfm:avm_writedata -> fpga_mem_inst:mrx_writedata
	wire   [25:0] fpga_mem_inst_mrx_bfm_m0_address;                                       // fpga_mem_inst_mrx_bfm:avm_address -> fpga_mem_inst:mrx_address
	wire          fpga_mem_inst_mrx_bfm_m0_write;                                         // fpga_mem_inst_mrx_bfm:avm_write -> fpga_mem_inst:mrx_write
	wire          fpga_mem_inst_mrx_bfm_m0_read;                                          // fpga_mem_inst_mrx_bfm:avm_read -> fpga_mem_inst:mrx_read
	wire  [127:0] fpga_mem_inst_mrx_bfm_m0_readdata;                                      // fpga_mem_inst:mrx_readdata -> fpga_mem_inst_mrx_bfm:avm_readdata
	wire          fpga_mem_inst_mrx_bfm_m0_debugaccess;                                   // fpga_mem_inst_mrx_bfm:avm_debugaccess -> fpga_mem_inst:mrx_debugaccess
	wire          fpga_mem_inst_mrx_bfm_m0_readdatavalid;                                 // fpga_mem_inst:mrx_readdatavalid -> fpga_mem_inst_mrx_bfm:avm_readdatavalid
	wire   [15:0] fpga_mem_inst_mrx_bfm_m0_byteenable;                                    // fpga_mem_inst_mrx_bfm:avm_byteenable -> fpga_mem_inst:mrx_byteenable
	wire          fpga_mem_inst_mr0_bfm_m0_waitrequest;                                   // fpga_mem_inst:mr0_waitrequest -> fpga_mem_inst_mr0_bfm:avm_waitrequest
	wire    [5:0] fpga_mem_inst_mr0_bfm_m0_burstcount;                                    // fpga_mem_inst_mr0_bfm:avm_burstcount -> fpga_mem_inst:mr0_burstcount
	wire  [127:0] fpga_mem_inst_mr0_bfm_m0_writedata;                                     // fpga_mem_inst_mr0_bfm:avm_writedata -> fpga_mem_inst:mr0_writedata
	wire   [25:0] fpga_mem_inst_mr0_bfm_m0_address;                                       // fpga_mem_inst_mr0_bfm:avm_address -> fpga_mem_inst:mr0_address
	wire          fpga_mem_inst_mr0_bfm_m0_write;                                         // fpga_mem_inst_mr0_bfm:avm_write -> fpga_mem_inst:mr0_write
	wire          fpga_mem_inst_mr0_bfm_m0_read;                                          // fpga_mem_inst_mr0_bfm:avm_read -> fpga_mem_inst:mr0_read
	wire  [127:0] fpga_mem_inst_mr0_bfm_m0_readdata;                                      // fpga_mem_inst:mr0_readdata -> fpga_mem_inst_mr0_bfm:avm_readdata
	wire          fpga_mem_inst_mr0_bfm_m0_debugaccess;                                   // fpga_mem_inst_mr0_bfm:avm_debugaccess -> fpga_mem_inst:mr0_debugaccess
	wire          fpga_mem_inst_mr0_bfm_m0_readdatavalid;                                 // fpga_mem_inst:mr0_readdatavalid -> fpga_mem_inst_mr0_bfm:avm_readdatavalid
	wire   [15:0] fpga_mem_inst_mr0_bfm_m0_byteenable;                                    // fpga_mem_inst_mr0_bfm:avm_byteenable -> fpga_mem_inst:mr0_byteenable
	wire          fpga_mem_inst_mr1_bfm_m0_waitrequest;                                   // fpga_mem_inst:mr1_waitrequest -> fpga_mem_inst_mr1_bfm:avm_waitrequest
	wire    [5:0] fpga_mem_inst_mr1_bfm_m0_burstcount;                                    // fpga_mem_inst_mr1_bfm:avm_burstcount -> fpga_mem_inst:mr1_burstcount
	wire  [127:0] fpga_mem_inst_mr1_bfm_m0_writedata;                                     // fpga_mem_inst_mr1_bfm:avm_writedata -> fpga_mem_inst:mr1_writedata
	wire   [25:0] fpga_mem_inst_mr1_bfm_m0_address;                                       // fpga_mem_inst_mr1_bfm:avm_address -> fpga_mem_inst:mr1_address
	wire          fpga_mem_inst_mr1_bfm_m0_write;                                         // fpga_mem_inst_mr1_bfm:avm_write -> fpga_mem_inst:mr1_write
	wire          fpga_mem_inst_mr1_bfm_m0_read;                                          // fpga_mem_inst_mr1_bfm:avm_read -> fpga_mem_inst:mr1_read
	wire  [127:0] fpga_mem_inst_mr1_bfm_m0_readdata;                                      // fpga_mem_inst:mr1_readdata -> fpga_mem_inst_mr1_bfm:avm_readdata
	wire          fpga_mem_inst_mr1_bfm_m0_debugaccess;                                   // fpga_mem_inst_mr1_bfm:avm_debugaccess -> fpga_mem_inst:mr1_debugaccess
	wire          fpga_mem_inst_mr1_bfm_m0_readdatavalid;                                 // fpga_mem_inst:mr1_readdatavalid -> fpga_mem_inst_mr1_bfm:avm_readdatavalid
	wire   [15:0] fpga_mem_inst_mr1_bfm_m0_byteenable;                                    // fpga_mem_inst_mr1_bfm:avm_byteenable -> fpga_mem_inst:mr1_byteenable
	wire          fpga_mem_inst_mr2_bfm_m0_waitrequest;                                   // fpga_mem_inst:mr2_waitrequest -> fpga_mem_inst_mr2_bfm:avm_waitrequest
	wire    [5:0] fpga_mem_inst_mr2_bfm_m0_burstcount;                                    // fpga_mem_inst_mr2_bfm:avm_burstcount -> fpga_mem_inst:mr2_burstcount
	wire  [127:0] fpga_mem_inst_mr2_bfm_m0_writedata;                                     // fpga_mem_inst_mr2_bfm:avm_writedata -> fpga_mem_inst:mr2_writedata
	wire   [25:0] fpga_mem_inst_mr2_bfm_m0_address;                                       // fpga_mem_inst_mr2_bfm:avm_address -> fpga_mem_inst:mr2_address
	wire          fpga_mem_inst_mr2_bfm_m0_write;                                         // fpga_mem_inst_mr2_bfm:avm_write -> fpga_mem_inst:mr2_write
	wire          fpga_mem_inst_mr2_bfm_m0_read;                                          // fpga_mem_inst_mr2_bfm:avm_read -> fpga_mem_inst:mr2_read
	wire  [127:0] fpga_mem_inst_mr2_bfm_m0_readdata;                                      // fpga_mem_inst:mr2_readdata -> fpga_mem_inst_mr2_bfm:avm_readdata
	wire          fpga_mem_inst_mr2_bfm_m0_debugaccess;                                   // fpga_mem_inst_mr2_bfm:avm_debugaccess -> fpga_mem_inst:mr2_debugaccess
	wire          fpga_mem_inst_mr2_bfm_m0_readdatavalid;                                 // fpga_mem_inst:mr2_readdatavalid -> fpga_mem_inst_mr2_bfm:avm_readdatavalid
	wire   [15:0] fpga_mem_inst_mr2_bfm_m0_byteenable;                                    // fpga_mem_inst_mr2_bfm:avm_byteenable -> fpga_mem_inst:mr2_byteenable
	wire          fpga_mem_inst_mr3_bfm_m0_waitrequest;                                   // fpga_mem_inst:mr3_waitrequest -> fpga_mem_inst_mr3_bfm:avm_waitrequest
	wire    [5:0] fpga_mem_inst_mr3_bfm_m0_burstcount;                                    // fpga_mem_inst_mr3_bfm:avm_burstcount -> fpga_mem_inst:mr3_burstcount
	wire  [127:0] fpga_mem_inst_mr3_bfm_m0_writedata;                                     // fpga_mem_inst_mr3_bfm:avm_writedata -> fpga_mem_inst:mr3_writedata
	wire   [25:0] fpga_mem_inst_mr3_bfm_m0_address;                                       // fpga_mem_inst_mr3_bfm:avm_address -> fpga_mem_inst:mr3_address
	wire          fpga_mem_inst_mr3_bfm_m0_write;                                         // fpga_mem_inst_mr3_bfm:avm_write -> fpga_mem_inst:mr3_write
	wire          fpga_mem_inst_mr3_bfm_m0_read;                                          // fpga_mem_inst_mr3_bfm:avm_read -> fpga_mem_inst:mr3_read
	wire  [127:0] fpga_mem_inst_mr3_bfm_m0_readdata;                                      // fpga_mem_inst:mr3_readdata -> fpga_mem_inst_mr3_bfm:avm_readdata
	wire          fpga_mem_inst_mr3_bfm_m0_debugaccess;                                   // fpga_mem_inst_mr3_bfm:avm_debugaccess -> fpga_mem_inst:mr3_debugaccess
	wire          fpga_mem_inst_mr3_bfm_m0_readdatavalid;                                 // fpga_mem_inst:mr3_readdatavalid -> fpga_mem_inst_mr3_bfm:avm_readdatavalid
	wire   [15:0] fpga_mem_inst_mr3_bfm_m0_byteenable;                                    // fpga_mem_inst_mr3_bfm:avm_byteenable -> fpga_mem_inst:mr3_byteenable
	wire          fpga_mem_inst_mwx_bfm_m0_waitrequest;                                   // fpga_mem_inst:mwx_waitrequest -> fpga_mem_inst_mwx_bfm:avm_waitrequest
	wire    [5:0] fpga_mem_inst_mwx_bfm_m0_burstcount;                                    // fpga_mem_inst_mwx_bfm:avm_burstcount -> fpga_mem_inst:mwx_burstcount
	wire  [127:0] fpga_mem_inst_mwx_bfm_m0_writedata;                                     // fpga_mem_inst_mwx_bfm:avm_writedata -> fpga_mem_inst:mwx_writedata
	wire   [25:0] fpga_mem_inst_mwx_bfm_m0_address;                                       // fpga_mem_inst_mwx_bfm:avm_address -> fpga_mem_inst:mwx_address
	wire          fpga_mem_inst_mwx_bfm_m0_write;                                         // fpga_mem_inst_mwx_bfm:avm_write -> fpga_mem_inst:mwx_write
	wire          fpga_mem_inst_mwx_bfm_m0_read;                                          // fpga_mem_inst_mwx_bfm:avm_read -> fpga_mem_inst:mwx_read
	wire  [127:0] fpga_mem_inst_mwx_bfm_m0_readdata;                                      // fpga_mem_inst:mwx_readdata -> fpga_mem_inst_mwx_bfm:avm_readdata
	wire          fpga_mem_inst_mwx_bfm_m0_debugaccess;                                   // fpga_mem_inst_mwx_bfm:avm_debugaccess -> fpga_mem_inst:mwx_debugaccess
	wire          fpga_mem_inst_mwx_bfm_m0_readdatavalid;                                 // fpga_mem_inst:mwx_readdatavalid -> fpga_mem_inst_mwx_bfm:avm_readdatavalid
	wire   [15:0] fpga_mem_inst_mwx_bfm_m0_byteenable;                                    // fpga_mem_inst_mwx_bfm:avm_byteenable -> fpga_mem_inst:mwx_byteenable
	wire          fpga_mem_inst_mw0_bfm_m0_waitrequest;                                   // fpga_mem_inst:mw0_waitrequest -> fpga_mem_inst_mw0_bfm:avm_waitrequest
	wire    [5:0] fpga_mem_inst_mw0_bfm_m0_burstcount;                                    // fpga_mem_inst_mw0_bfm:avm_burstcount -> fpga_mem_inst:mw0_burstcount
	wire  [127:0] fpga_mem_inst_mw0_bfm_m0_writedata;                                     // fpga_mem_inst_mw0_bfm:avm_writedata -> fpga_mem_inst:mw0_writedata
	wire   [25:0] fpga_mem_inst_mw0_bfm_m0_address;                                       // fpga_mem_inst_mw0_bfm:avm_address -> fpga_mem_inst:mw0_address
	wire          fpga_mem_inst_mw0_bfm_m0_write;                                         // fpga_mem_inst_mw0_bfm:avm_write -> fpga_mem_inst:mw0_write
	wire          fpga_mem_inst_mw0_bfm_m0_read;                                          // fpga_mem_inst_mw0_bfm:avm_read -> fpga_mem_inst:mw0_read
	wire  [127:0] fpga_mem_inst_mw0_bfm_m0_readdata;                                      // fpga_mem_inst:mw0_readdata -> fpga_mem_inst_mw0_bfm:avm_readdata
	wire          fpga_mem_inst_mw0_bfm_m0_debugaccess;                                   // fpga_mem_inst_mw0_bfm:avm_debugaccess -> fpga_mem_inst:mw0_debugaccess
	wire          fpga_mem_inst_mw0_bfm_m0_readdatavalid;                                 // fpga_mem_inst:mw0_readdatavalid -> fpga_mem_inst_mw0_bfm:avm_readdatavalid
	wire   [15:0] fpga_mem_inst_mw0_bfm_m0_byteenable;                                    // fpga_mem_inst_mw0_bfm:avm_byteenable -> fpga_mem_inst:mw0_byteenable
	wire          fpga_mem_inst_mw1_bfm_m0_waitrequest;                                   // fpga_mem_inst:mw1_waitrequest -> fpga_mem_inst_mw1_bfm:avm_waitrequest
	wire    [5:0] fpga_mem_inst_mw1_bfm_m0_burstcount;                                    // fpga_mem_inst_mw1_bfm:avm_burstcount -> fpga_mem_inst:mw1_burstcount
	wire  [127:0] fpga_mem_inst_mw1_bfm_m0_writedata;                                     // fpga_mem_inst_mw1_bfm:avm_writedata -> fpga_mem_inst:mw1_writedata
	wire   [25:0] fpga_mem_inst_mw1_bfm_m0_address;                                       // fpga_mem_inst_mw1_bfm:avm_address -> fpga_mem_inst:mw1_address
	wire          fpga_mem_inst_mw1_bfm_m0_write;                                         // fpga_mem_inst_mw1_bfm:avm_write -> fpga_mem_inst:mw1_write
	wire          fpga_mem_inst_mw1_bfm_m0_read;                                          // fpga_mem_inst_mw1_bfm:avm_read -> fpga_mem_inst:mw1_read
	wire  [127:0] fpga_mem_inst_mw1_bfm_m0_readdata;                                      // fpga_mem_inst:mw1_readdata -> fpga_mem_inst_mw1_bfm:avm_readdata
	wire          fpga_mem_inst_mw1_bfm_m0_debugaccess;                                   // fpga_mem_inst_mw1_bfm:avm_debugaccess -> fpga_mem_inst:mw1_debugaccess
	wire          fpga_mem_inst_mw1_bfm_m0_readdatavalid;                                 // fpga_mem_inst:mw1_readdatavalid -> fpga_mem_inst_mw1_bfm:avm_readdatavalid
	wire   [15:0] fpga_mem_inst_mw1_bfm_m0_byteenable;                                    // fpga_mem_inst_mw1_bfm:avm_byteenable -> fpga_mem_inst:mw1_byteenable
	wire          fpga_mem_inst_mw2_bfm_m0_waitrequest;                                   // fpga_mem_inst:mw2_waitrequest -> fpga_mem_inst_mw2_bfm:avm_waitrequest
	wire    [5:0] fpga_mem_inst_mw2_bfm_m0_burstcount;                                    // fpga_mem_inst_mw2_bfm:avm_burstcount -> fpga_mem_inst:mw2_burstcount
	wire  [127:0] fpga_mem_inst_mw2_bfm_m0_writedata;                                     // fpga_mem_inst_mw2_bfm:avm_writedata -> fpga_mem_inst:mw2_writedata
	wire   [25:0] fpga_mem_inst_mw2_bfm_m0_address;                                       // fpga_mem_inst_mw2_bfm:avm_address -> fpga_mem_inst:mw2_address
	wire          fpga_mem_inst_mw2_bfm_m0_write;                                         // fpga_mem_inst_mw2_bfm:avm_write -> fpga_mem_inst:mw2_write
	wire          fpga_mem_inst_mw2_bfm_m0_read;                                          // fpga_mem_inst_mw2_bfm:avm_read -> fpga_mem_inst:mw2_read
	wire  [127:0] fpga_mem_inst_mw2_bfm_m0_readdata;                                      // fpga_mem_inst:mw2_readdata -> fpga_mem_inst_mw2_bfm:avm_readdata
	wire          fpga_mem_inst_mw2_bfm_m0_debugaccess;                                   // fpga_mem_inst_mw2_bfm:avm_debugaccess -> fpga_mem_inst:mw2_debugaccess
	wire          fpga_mem_inst_mw2_bfm_m0_readdatavalid;                                 // fpga_mem_inst:mw2_readdatavalid -> fpga_mem_inst_mw2_bfm:avm_readdatavalid
	wire   [15:0] fpga_mem_inst_mw2_bfm_m0_byteenable;                                    // fpga_mem_inst_mw2_bfm:avm_byteenable -> fpga_mem_inst:mw2_byteenable
	wire          fpga_mem_inst_mw3_bfm_m0_waitrequest;                                   // fpga_mem_inst:mw3_waitrequest -> fpga_mem_inst_mw3_bfm:avm_waitrequest
	wire    [5:0] fpga_mem_inst_mw3_bfm_m0_burstcount;                                    // fpga_mem_inst_mw3_bfm:avm_burstcount -> fpga_mem_inst:mw3_burstcount
	wire  [127:0] fpga_mem_inst_mw3_bfm_m0_writedata;                                     // fpga_mem_inst_mw3_bfm:avm_writedata -> fpga_mem_inst:mw3_writedata
	wire   [25:0] fpga_mem_inst_mw3_bfm_m0_address;                                       // fpga_mem_inst_mw3_bfm:avm_address -> fpga_mem_inst:mw3_address
	wire          fpga_mem_inst_mw3_bfm_m0_write;                                         // fpga_mem_inst_mw3_bfm:avm_write -> fpga_mem_inst:mw3_write
	wire          fpga_mem_inst_mw3_bfm_m0_read;                                          // fpga_mem_inst_mw3_bfm:avm_read -> fpga_mem_inst:mw3_read
	wire  [127:0] fpga_mem_inst_mw3_bfm_m0_readdata;                                      // fpga_mem_inst:mw3_readdata -> fpga_mem_inst_mw3_bfm:avm_readdata
	wire          fpga_mem_inst_mw3_bfm_m0_debugaccess;                                   // fpga_mem_inst_mw3_bfm:avm_debugaccess -> fpga_mem_inst:mw3_debugaccess
	wire          fpga_mem_inst_mw3_bfm_m0_readdatavalid;                                 // fpga_mem_inst:mw3_readdatavalid -> fpga_mem_inst_mw3_bfm:avm_readdatavalid
	wire   [15:0] fpga_mem_inst_mw3_bfm_m0_byteenable;                                    // fpga_mem_inst_mw3_bfm:avm_byteenable -> fpga_mem_inst:mw3_byteenable
	wire          fpga_mem_inst_hps_bfm_m0_waitrequest;                                   // fpga_mem_inst:hps_waitrequest -> fpga_mem_inst_hps_bfm:avm_waitrequest
	wire    [5:0] fpga_mem_inst_hps_bfm_m0_burstcount;                                    // fpga_mem_inst_hps_bfm:avm_burstcount -> fpga_mem_inst:hps_burstcount
	wire  [127:0] fpga_mem_inst_hps_bfm_m0_writedata;                                     // fpga_mem_inst_hps_bfm:avm_writedata -> fpga_mem_inst:hps_writedata
	wire   [25:0] fpga_mem_inst_hps_bfm_m0_address;                                       // fpga_mem_inst_hps_bfm:avm_address -> fpga_mem_inst:hps_address
	wire          fpga_mem_inst_hps_bfm_m0_write;                                         // fpga_mem_inst_hps_bfm:avm_write -> fpga_mem_inst:hps_write
	wire          fpga_mem_inst_hps_bfm_m0_read;                                          // fpga_mem_inst_hps_bfm:avm_read -> fpga_mem_inst:hps_read
	wire  [127:0] fpga_mem_inst_hps_bfm_m0_readdata;                                      // fpga_mem_inst:hps_readdata -> fpga_mem_inst_hps_bfm:avm_readdata
	wire          fpga_mem_inst_hps_bfm_m0_debugaccess;                                   // fpga_mem_inst_hps_bfm:avm_debugaccess -> fpga_mem_inst:hps_debugaccess
	wire          fpga_mem_inst_hps_bfm_m0_readdatavalid;                                 // fpga_mem_inst:hps_readdatavalid -> fpga_mem_inst_hps_bfm:avm_readdatavalid
	wire   [15:0] fpga_mem_inst_hps_bfm_m0_byteenable;                                    // fpga_mem_inst_hps_bfm:avm_byteenable -> fpga_mem_inst:hps_byteenable
	wire    [0:0] fpga_mem_inst_memory_0_mem_odt;                                         // fpga_mem_inst:memory_0_mem_odt -> mem_if_ddr3_emif_0_mem_model:mem_odt
	wire    [0:0] fpga_mem_inst_memory_0_mem_cs_n;                                        // fpga_mem_inst:memory_0_mem_cs_n -> mem_if_ddr3_emif_0_mem_model:mem_cs_n
	wire   [14:0] fpga_mem_inst_memory_0_mem_a;                                           // fpga_mem_inst:memory_0_mem_a -> mem_if_ddr3_emif_0_mem_model:mem_a
	wire    [0:0] fpga_mem_inst_memory_0_mem_ck_n;                                        // fpga_mem_inst:memory_0_mem_ck_n -> mem_if_ddr3_emif_0_mem_model:mem_ck_n
	wire    [0:0] fpga_mem_inst_memory_0_mem_ras_n;                                       // fpga_mem_inst:memory_0_mem_ras_n -> mem_if_ddr3_emif_0_mem_model:mem_ras_n
	wire    [0:0] fpga_mem_inst_memory_0_mem_cke;                                         // fpga_mem_inst:memory_0_mem_cke -> mem_if_ddr3_emif_0_mem_model:mem_cke
	wire    [3:0] fpga_mem_inst_memory_0_mem_dqs;                                         // [] -> [fpga_mem_inst:memory_0_mem_dqs, mem_if_ddr3_emif_0_mem_model:mem_dqs]
	wire    [0:0] fpga_mem_inst_memory_0_mem_we_n;                                        // fpga_mem_inst:memory_0_mem_we_n -> mem_if_ddr3_emif_0_mem_model:mem_we_n
	wire    [2:0] fpga_mem_inst_memory_0_mem_ba;                                          // fpga_mem_inst:memory_0_mem_ba -> mem_if_ddr3_emif_0_mem_model:mem_ba
	wire   [31:0] fpga_mem_inst_memory_0_mem_dq;                                          // [] -> [fpga_mem_inst:memory_0_mem_dq, mem_if_ddr3_emif_0_mem_model:mem_dq]
	wire    [0:0] fpga_mem_inst_memory_0_mem_ck;                                          // fpga_mem_inst:memory_0_mem_ck -> mem_if_ddr3_emif_0_mem_model:mem_ck
	wire          fpga_mem_inst_memory_0_mem_reset_n;                                     // fpga_mem_inst:memory_0_mem_reset_n -> mem_if_ddr3_emif_0_mem_model:mem_reset_n
	wire    [3:0] fpga_mem_inst_memory_0_mem_dm;                                          // fpga_mem_inst:memory_0_mem_dm -> mem_if_ddr3_emif_0_mem_model:mem_dm
	wire    [0:0] fpga_mem_inst_memory_0_mem_cas_n;                                       // fpga_mem_inst:memory_0_mem_cas_n -> mem_if_ddr3_emif_0_mem_model:mem_cas_n
	wire    [3:0] fpga_mem_inst_memory_0_mem_dqs_n;                                       // [] -> [fpga_mem_inst:memory_0_mem_dqs_n, mem_if_ddr3_emif_0_mem_model:mem_dqs_n]
	wire          rst_controller_reset_out_reset;                                         // rst_controller:reset_out -> [fpga_mem_inst_hps_bfm:reset, fpga_mem_inst_mr0_bfm:reset, fpga_mem_inst_mr1_bfm:reset, fpga_mem_inst_mr2_bfm:reset, fpga_mem_inst_mr3_bfm:reset, fpga_mem_inst_mrx_bfm:reset, fpga_mem_inst_mw0_bfm:reset, fpga_mem_inst_mw1_bfm:reset, fpga_mem_inst_mw2_bfm:reset, fpga_mem_inst_mw3_bfm:reset, fpga_mem_inst_mwx_bfm:reset]

	fpga_mem fpga_mem_inst (
		.clk_clk                                                  (fpga_mem_inst_clk_bfm_clk_clk),                                          //                            clk.clk
		.reset_reset_n                                            (fpga_mem_inst_reset_bfm_reset_reset),                                    //                          reset.reset_n
		.memory_0_mem_a                                           (fpga_mem_inst_memory_0_mem_a),                                           //                       memory_0.mem_a
		.memory_0_mem_ba                                          (fpga_mem_inst_memory_0_mem_ba),                                          //                               .mem_ba
		.memory_0_mem_ck                                          (fpga_mem_inst_memory_0_mem_ck),                                          //                               .mem_ck
		.memory_0_mem_ck_n                                        (fpga_mem_inst_memory_0_mem_ck_n),                                        //                               .mem_ck_n
		.memory_0_mem_cke                                         (fpga_mem_inst_memory_0_mem_cke),                                         //                               .mem_cke
		.memory_0_mem_cs_n                                        (fpga_mem_inst_memory_0_mem_cs_n),                                        //                               .mem_cs_n
		.memory_0_mem_dm                                          (fpga_mem_inst_memory_0_mem_dm),                                          //                               .mem_dm
		.memory_0_mem_ras_n                                       (fpga_mem_inst_memory_0_mem_ras_n),                                       //                               .mem_ras_n
		.memory_0_mem_cas_n                                       (fpga_mem_inst_memory_0_mem_cas_n),                                       //                               .mem_cas_n
		.memory_0_mem_we_n                                        (fpga_mem_inst_memory_0_mem_we_n),                                        //                               .mem_we_n
		.memory_0_mem_reset_n                                     (fpga_mem_inst_memory_0_mem_reset_n),                                     //                               .mem_reset_n
		.memory_0_mem_dq                                          (fpga_mem_inst_memory_0_mem_dq),                                          //                               .mem_dq
		.memory_0_mem_dqs                                         (fpga_mem_inst_memory_0_mem_dqs),                                         //                               .mem_dqs
		.memory_0_mem_dqs_n                                       (fpga_mem_inst_memory_0_mem_dqs_n),                                       //                               .mem_dqs_n
		.memory_0_mem_odt                                         (fpga_mem_inst_memory_0_mem_odt),                                         //                               .mem_odt
		.oct_rzqin                                                (fpga_mem_inst_oct_bfm_conduit_rzqin),                                    //                            oct.rzqin
		.mem_if_ddr3_emif_0_status_local_init_done                (fpga_mem_inst_mem_if_ddr3_emif_0_status_local_init_done),                //      mem_if_ddr3_emif_0_status.local_init_done
		.mem_if_ddr3_emif_0_status_local_cal_success              (fpga_mem_inst_mem_if_ddr3_emif_0_status_local_cal_success),              //                               .local_cal_success
		.mem_if_ddr3_emif_0_status_local_cal_fail                 (fpga_mem_inst_mem_if_ddr3_emif_0_status_local_cal_fail),                 //                               .local_cal_fail
		.mem_if_ddr3_emif_0_pll_sharing_pll_mem_clk               (fpga_mem_inst_mem_if_ddr3_emif_0_pll_sharing_pll_mem_clk),               // mem_if_ddr3_emif_0_pll_sharing.pll_mem_clk
		.mem_if_ddr3_emif_0_pll_sharing_pll_write_clk             (fpga_mem_inst_mem_if_ddr3_emif_0_pll_sharing_pll_write_clk),             //                               .pll_write_clk
		.mem_if_ddr3_emif_0_pll_sharing_pll_locked                (fpga_mem_inst_mem_if_ddr3_emif_0_pll_sharing_pll_locked),                //                               .pll_locked
		.mem_if_ddr3_emif_0_pll_sharing_pll_write_clk_pre_phy_clk (fpga_mem_inst_mem_if_ddr3_emif_0_pll_sharing_pll_write_clk_pre_phy_clk), //                               .pll_write_clk_pre_phy_clk
		.mem_if_ddr3_emif_0_pll_sharing_pll_addr_cmd_clk          (fpga_mem_inst_mem_if_ddr3_emif_0_pll_sharing_pll_addr_cmd_clk),          //                               .pll_addr_cmd_clk
		.mem_if_ddr3_emif_0_pll_sharing_pll_avl_clk               (fpga_mem_inst_mem_if_ddr3_emif_0_pll_sharing_pll_avl_clk),               //                               .pll_avl_clk
		.mem_if_ddr3_emif_0_pll_sharing_pll_config_clk            (fpga_mem_inst_mem_if_ddr3_emif_0_pll_sharing_pll_config_clk),            //                               .pll_config_clk
		.mem_if_ddr3_emif_0_pll_sharing_pll_dr_clk                (fpga_mem_inst_mem_if_ddr3_emif_0_pll_sharing_pll_dr_clk),                //                               .pll_dr_clk
		.mem_if_ddr3_emif_0_pll_sharing_pll_dr_clk_pre_phy_clk    (fpga_mem_inst_mem_if_ddr3_emif_0_pll_sharing_pll_dr_clk_pre_phy_clk),    //                               .pll_dr_clk_pre_phy_clk
		.mem_if_ddr3_emif_0_pll_sharing_pll_mem_phy_clk           (fpga_mem_inst_mem_if_ddr3_emif_0_pll_sharing_pll_mem_phy_clk),           //                               .pll_mem_phy_clk
		.mem_if_ddr3_emif_0_pll_sharing_afi_phy_clk               (fpga_mem_inst_mem_if_ddr3_emif_0_pll_sharing_afi_phy_clk),               //                               .afi_phy_clk
		.mem_if_ddr3_emif_0_pll_sharing_pll_avl_phy_clk           (fpga_mem_inst_mem_if_ddr3_emif_0_pll_sharing_pll_avl_phy_clk),           //                               .pll_avl_phy_clk
		.afi_clk_clk                                              (fpga_mem_inst_afi_clk_clk),                                              //                        afi_clk.clk
		.mrx_waitrequest                                          (fpga_mem_inst_mrx_bfm_m0_waitrequest),                                   //                            mrx.waitrequest
		.mrx_readdata                                             (fpga_mem_inst_mrx_bfm_m0_readdata),                                      //                               .readdata
		.mrx_readdatavalid                                        (fpga_mem_inst_mrx_bfm_m0_readdatavalid),                                 //                               .readdatavalid
		.mrx_burstcount                                           (fpga_mem_inst_mrx_bfm_m0_burstcount),                                    //                               .burstcount
		.mrx_writedata                                            (fpga_mem_inst_mrx_bfm_m0_writedata),                                     //                               .writedata
		.mrx_address                                              (fpga_mem_inst_mrx_bfm_m0_address),                                       //                               .address
		.mrx_write                                                (fpga_mem_inst_mrx_bfm_m0_write),                                         //                               .write
		.mrx_read                                                 (fpga_mem_inst_mrx_bfm_m0_read),                                          //                               .read
		.mrx_byteenable                                           (fpga_mem_inst_mrx_bfm_m0_byteenable),                                    //                               .byteenable
		.mrx_debugaccess                                          (fpga_mem_inst_mrx_bfm_m0_debugaccess),                                   //                               .debugaccess
		.mr0_waitrequest                                          (fpga_mem_inst_mr0_bfm_m0_waitrequest),                                   //                            mr0.waitrequest
		.mr0_readdata                                             (fpga_mem_inst_mr0_bfm_m0_readdata),                                      //                               .readdata
		.mr0_readdatavalid                                        (fpga_mem_inst_mr0_bfm_m0_readdatavalid),                                 //                               .readdatavalid
		.mr0_burstcount                                           (fpga_mem_inst_mr0_bfm_m0_burstcount),                                    //                               .burstcount
		.mr0_writedata                                            (fpga_mem_inst_mr0_bfm_m0_writedata),                                     //                               .writedata
		.mr0_address                                              (fpga_mem_inst_mr0_bfm_m0_address),                                       //                               .address
		.mr0_write                                                (fpga_mem_inst_mr0_bfm_m0_write),                                         //                               .write
		.mr0_read                                                 (fpga_mem_inst_mr0_bfm_m0_read),                                          //                               .read
		.mr0_byteenable                                           (fpga_mem_inst_mr0_bfm_m0_byteenable),                                    //                               .byteenable
		.mr0_debugaccess                                          (fpga_mem_inst_mr0_bfm_m0_debugaccess),                                   //                               .debugaccess
		.mr1_waitrequest                                          (fpga_mem_inst_mr1_bfm_m0_waitrequest),                                   //                            mr1.waitrequest
		.mr1_readdata                                             (fpga_mem_inst_mr1_bfm_m0_readdata),                                      //                               .readdata
		.mr1_readdatavalid                                        (fpga_mem_inst_mr1_bfm_m0_readdatavalid),                                 //                               .readdatavalid
		.mr1_burstcount                                           (fpga_mem_inst_mr1_bfm_m0_burstcount),                                    //                               .burstcount
		.mr1_writedata                                            (fpga_mem_inst_mr1_bfm_m0_writedata),                                     //                               .writedata
		.mr1_address                                              (fpga_mem_inst_mr1_bfm_m0_address),                                       //                               .address
		.mr1_write                                                (fpga_mem_inst_mr1_bfm_m0_write),                                         //                               .write
		.mr1_read                                                 (fpga_mem_inst_mr1_bfm_m0_read),                                          //                               .read
		.mr1_byteenable                                           (fpga_mem_inst_mr1_bfm_m0_byteenable),                                    //                               .byteenable
		.mr1_debugaccess                                          (fpga_mem_inst_mr1_bfm_m0_debugaccess),                                   //                               .debugaccess
		.mr2_waitrequest                                          (fpga_mem_inst_mr2_bfm_m0_waitrequest),                                   //                            mr2.waitrequest
		.mr2_readdata                                             (fpga_mem_inst_mr2_bfm_m0_readdata),                                      //                               .readdata
		.mr2_readdatavalid                                        (fpga_mem_inst_mr2_bfm_m0_readdatavalid),                                 //                               .readdatavalid
		.mr2_burstcount                                           (fpga_mem_inst_mr2_bfm_m0_burstcount),                                    //                               .burstcount
		.mr2_writedata                                            (fpga_mem_inst_mr2_bfm_m0_writedata),                                     //                               .writedata
		.mr2_address                                              (fpga_mem_inst_mr2_bfm_m0_address),                                       //                               .address
		.mr2_write                                                (fpga_mem_inst_mr2_bfm_m0_write),                                         //                               .write
		.mr2_read                                                 (fpga_mem_inst_mr2_bfm_m0_read),                                          //                               .read
		.mr2_byteenable                                           (fpga_mem_inst_mr2_bfm_m0_byteenable),                                    //                               .byteenable
		.mr2_debugaccess                                          (fpga_mem_inst_mr2_bfm_m0_debugaccess),                                   //                               .debugaccess
		.mr3_waitrequest                                          (fpga_mem_inst_mr3_bfm_m0_waitrequest),                                   //                            mr3.waitrequest
		.mr3_readdata                                             (fpga_mem_inst_mr3_bfm_m0_readdata),                                      //                               .readdata
		.mr3_readdatavalid                                        (fpga_mem_inst_mr3_bfm_m0_readdatavalid),                                 //                               .readdatavalid
		.mr3_burstcount                                           (fpga_mem_inst_mr3_bfm_m0_burstcount),                                    //                               .burstcount
		.mr3_writedata                                            (fpga_mem_inst_mr3_bfm_m0_writedata),                                     //                               .writedata
		.mr3_address                                              (fpga_mem_inst_mr3_bfm_m0_address),                                       //                               .address
		.mr3_write                                                (fpga_mem_inst_mr3_bfm_m0_write),                                         //                               .write
		.mr3_read                                                 (fpga_mem_inst_mr3_bfm_m0_read),                                          //                               .read
		.mr3_byteenable                                           (fpga_mem_inst_mr3_bfm_m0_byteenable),                                    //                               .byteenable
		.mr3_debugaccess                                          (fpga_mem_inst_mr3_bfm_m0_debugaccess),                                   //                               .debugaccess
		.mwx_waitrequest                                          (fpga_mem_inst_mwx_bfm_m0_waitrequest),                                   //                            mwx.waitrequest
		.mwx_readdata                                             (fpga_mem_inst_mwx_bfm_m0_readdata),                                      //                               .readdata
		.mwx_readdatavalid                                        (fpga_mem_inst_mwx_bfm_m0_readdatavalid),                                 //                               .readdatavalid
		.mwx_burstcount                                           (fpga_mem_inst_mwx_bfm_m0_burstcount),                                    //                               .burstcount
		.mwx_writedata                                            (fpga_mem_inst_mwx_bfm_m0_writedata),                                     //                               .writedata
		.mwx_address                                              (fpga_mem_inst_mwx_bfm_m0_address),                                       //                               .address
		.mwx_write                                                (fpga_mem_inst_mwx_bfm_m0_write),                                         //                               .write
		.mwx_read                                                 (fpga_mem_inst_mwx_bfm_m0_read),                                          //                               .read
		.mwx_byteenable                                           (fpga_mem_inst_mwx_bfm_m0_byteenable),                                    //                               .byteenable
		.mwx_debugaccess                                          (fpga_mem_inst_mwx_bfm_m0_debugaccess),                                   //                               .debugaccess
		.mw0_waitrequest                                          (fpga_mem_inst_mw0_bfm_m0_waitrequest),                                   //                            mw0.waitrequest
		.mw0_readdata                                             (fpga_mem_inst_mw0_bfm_m0_readdata),                                      //                               .readdata
		.mw0_readdatavalid                                        (fpga_mem_inst_mw0_bfm_m0_readdatavalid),                                 //                               .readdatavalid
		.mw0_burstcount                                           (fpga_mem_inst_mw0_bfm_m0_burstcount),                                    //                               .burstcount
		.mw0_writedata                                            (fpga_mem_inst_mw0_bfm_m0_writedata),                                     //                               .writedata
		.mw0_address                                              (fpga_mem_inst_mw0_bfm_m0_address),                                       //                               .address
		.mw0_write                                                (fpga_mem_inst_mw0_bfm_m0_write),                                         //                               .write
		.mw0_read                                                 (fpga_mem_inst_mw0_bfm_m0_read),                                          //                               .read
		.mw0_byteenable                                           (fpga_mem_inst_mw0_bfm_m0_byteenable),                                    //                               .byteenable
		.mw0_debugaccess                                          (fpga_mem_inst_mw0_bfm_m0_debugaccess),                                   //                               .debugaccess
		.mw1_waitrequest                                          (fpga_mem_inst_mw1_bfm_m0_waitrequest),                                   //                            mw1.waitrequest
		.mw1_readdata                                             (fpga_mem_inst_mw1_bfm_m0_readdata),                                      //                               .readdata
		.mw1_readdatavalid                                        (fpga_mem_inst_mw1_bfm_m0_readdatavalid),                                 //                               .readdatavalid
		.mw1_burstcount                                           (fpga_mem_inst_mw1_bfm_m0_burstcount),                                    //                               .burstcount
		.mw1_writedata                                            (fpga_mem_inst_mw1_bfm_m0_writedata),                                     //                               .writedata
		.mw1_address                                              (fpga_mem_inst_mw1_bfm_m0_address),                                       //                               .address
		.mw1_write                                                (fpga_mem_inst_mw1_bfm_m0_write),                                         //                               .write
		.mw1_read                                                 (fpga_mem_inst_mw1_bfm_m0_read),                                          //                               .read
		.mw1_byteenable                                           (fpga_mem_inst_mw1_bfm_m0_byteenable),                                    //                               .byteenable
		.mw1_debugaccess                                          (fpga_mem_inst_mw1_bfm_m0_debugaccess),                                   //                               .debugaccess
		.mw2_waitrequest                                          (fpga_mem_inst_mw2_bfm_m0_waitrequest),                                   //                            mw2.waitrequest
		.mw2_readdata                                             (fpga_mem_inst_mw2_bfm_m0_readdata),                                      //                               .readdata
		.mw2_readdatavalid                                        (fpga_mem_inst_mw2_bfm_m0_readdatavalid),                                 //                               .readdatavalid
		.mw2_burstcount                                           (fpga_mem_inst_mw2_bfm_m0_burstcount),                                    //                               .burstcount
		.mw2_writedata                                            (fpga_mem_inst_mw2_bfm_m0_writedata),                                     //                               .writedata
		.mw2_address                                              (fpga_mem_inst_mw2_bfm_m0_address),                                       //                               .address
		.mw2_write                                                (fpga_mem_inst_mw2_bfm_m0_write),                                         //                               .write
		.mw2_read                                                 (fpga_mem_inst_mw2_bfm_m0_read),                                          //                               .read
		.mw2_byteenable                                           (fpga_mem_inst_mw2_bfm_m0_byteenable),                                    //                               .byteenable
		.mw2_debugaccess                                          (fpga_mem_inst_mw2_bfm_m0_debugaccess),                                   //                               .debugaccess
		.mw3_waitrequest                                          (fpga_mem_inst_mw3_bfm_m0_waitrequest),                                   //                            mw3.waitrequest
		.mw3_readdata                                             (fpga_mem_inst_mw3_bfm_m0_readdata),                                      //                               .readdata
		.mw3_readdatavalid                                        (fpga_mem_inst_mw3_bfm_m0_readdatavalid),                                 //                               .readdatavalid
		.mw3_burstcount                                           (fpga_mem_inst_mw3_bfm_m0_burstcount),                                    //                               .burstcount
		.mw3_writedata                                            (fpga_mem_inst_mw3_bfm_m0_writedata),                                     //                               .writedata
		.mw3_address                                              (fpga_mem_inst_mw3_bfm_m0_address),                                       //                               .address
		.mw3_write                                                (fpga_mem_inst_mw3_bfm_m0_write),                                         //                               .write
		.mw3_read                                                 (fpga_mem_inst_mw3_bfm_m0_read),                                          //                               .read
		.mw3_byteenable                                           (fpga_mem_inst_mw3_bfm_m0_byteenable),                                    //                               .byteenable
		.mw3_debugaccess                                          (fpga_mem_inst_mw3_bfm_m0_debugaccess),                                   //                               .debugaccess
		.hps_waitrequest                                          (fpga_mem_inst_hps_bfm_m0_waitrequest),                                   //                            hps.waitrequest
		.hps_readdata                                             (fpga_mem_inst_hps_bfm_m0_readdata),                                      //                               .readdata
		.hps_readdatavalid                                        (fpga_mem_inst_hps_bfm_m0_readdatavalid),                                 //                               .readdatavalid
		.hps_burstcount                                           (fpga_mem_inst_hps_bfm_m0_burstcount),                                    //                               .burstcount
		.hps_writedata                                            (fpga_mem_inst_hps_bfm_m0_writedata),                                     //                               .writedata
		.hps_address                                              (fpga_mem_inst_hps_bfm_m0_address),                                       //                               .address
		.hps_write                                                (fpga_mem_inst_hps_bfm_m0_write),                                         //                               .write
		.hps_read                                                 (fpga_mem_inst_hps_bfm_m0_read),                                          //                               .read
		.hps_byteenable                                           (fpga_mem_inst_hps_bfm_m0_byteenable),                                    //                               .byteenable
		.hps_debugaccess                                          (fpga_mem_inst_hps_bfm_m0_debugaccess)                                    //                               .debugaccess
	);

	altera_avalon_clock_source #(
		.CLOCK_RATE (50000000),
		.CLOCK_UNIT (1)
	) fpga_mem_inst_clk_bfm (
		.clk (fpga_mem_inst_clk_bfm_clk_clk)  // clk.clk
	);

	altera_avalon_reset_source #(
		.ASSERT_HIGH_RESET    (0),
		.INITIAL_RESET_CYCLES (50)
	) fpga_mem_inst_reset_bfm (
		.reset (fpga_mem_inst_reset_bfm_reset_reset), // reset.reset_n
		.clk   (fpga_mem_inst_clk_bfm_clk_clk)        //   clk.clk
	);

	altera_conduit_bfm fpga_mem_inst_oct_bfm (
		.sig_rzqin (fpga_mem_inst_oct_bfm_conduit_rzqin)  // conduit.rzqin
	);

	altera_conduit_bfm_0002 fpga_mem_inst_mem_if_ddr3_emif_0_status_bfm (
		.sig_local_init_done   (fpga_mem_inst_mem_if_ddr3_emif_0_status_local_init_done),   // conduit.local_init_done
		.sig_local_cal_success (fpga_mem_inst_mem_if_ddr3_emif_0_status_local_cal_success), //        .local_cal_success
		.sig_local_cal_fail    (fpga_mem_inst_mem_if_ddr3_emif_0_status_local_cal_fail)     //        .local_cal_fail
	);

	altera_conduit_bfm_0003 fpga_mem_inst_mem_if_ddr3_emif_0_pll_sharing_bfm (
		.sig_pll_mem_clk               (fpga_mem_inst_mem_if_ddr3_emif_0_pll_sharing_pll_mem_clk),               // conduit.pll_mem_clk
		.sig_pll_write_clk             (fpga_mem_inst_mem_if_ddr3_emif_0_pll_sharing_pll_write_clk),             //        .pll_write_clk
		.sig_pll_locked                (fpga_mem_inst_mem_if_ddr3_emif_0_pll_sharing_pll_locked),                //        .pll_locked
		.sig_pll_write_clk_pre_phy_clk (fpga_mem_inst_mem_if_ddr3_emif_0_pll_sharing_pll_write_clk_pre_phy_clk), //        .pll_write_clk_pre_phy_clk
		.sig_pll_addr_cmd_clk          (fpga_mem_inst_mem_if_ddr3_emif_0_pll_sharing_pll_addr_cmd_clk),          //        .pll_addr_cmd_clk
		.sig_pll_avl_clk               (fpga_mem_inst_mem_if_ddr3_emif_0_pll_sharing_pll_avl_clk),               //        .pll_avl_clk
		.sig_pll_config_clk            (fpga_mem_inst_mem_if_ddr3_emif_0_pll_sharing_pll_config_clk),            //        .pll_config_clk
		.sig_pll_dr_clk                (fpga_mem_inst_mem_if_ddr3_emif_0_pll_sharing_pll_dr_clk),                //        .pll_dr_clk
		.sig_pll_dr_clk_pre_phy_clk    (fpga_mem_inst_mem_if_ddr3_emif_0_pll_sharing_pll_dr_clk_pre_phy_clk),    //        .pll_dr_clk_pre_phy_clk
		.sig_pll_mem_phy_clk           (fpga_mem_inst_mem_if_ddr3_emif_0_pll_sharing_pll_mem_phy_clk),           //        .pll_mem_phy_clk
		.sig_afi_phy_clk               (fpga_mem_inst_mem_if_ddr3_emif_0_pll_sharing_afi_phy_clk),               //        .afi_phy_clk
		.sig_pll_avl_phy_clk           (fpga_mem_inst_mem_if_ddr3_emif_0_pll_sharing_pll_avl_phy_clk)            //        .pll_avl_phy_clk
	);

	altera_avalon_mm_master_bfm #(
		.AV_ADDRESS_W               (26),
		.AV_SYMBOL_W                (8),
		.AV_NUMSYMBOLS              (16),
		.AV_BURSTCOUNT_W            (6),
		.AV_READRESPONSE_W          (1),
		.AV_WRITERESPONSE_W         (1),
		.USE_READ                   (1),
		.USE_WRITE                  (1),
		.USE_ADDRESS                (1),
		.USE_BYTE_ENABLE            (1),
		.USE_BURSTCOUNT             (1),
		.USE_READ_DATA              (1),
		.USE_READ_DATA_VALID        (1),
		.USE_WRITE_DATA             (1),
		.USE_BEGIN_TRANSFER         (0),
		.USE_BEGIN_BURST_TRANSFER   (0),
		.USE_WAIT_REQUEST           (1),
		.USE_TRANSACTIONID          (0),
		.USE_WRITERESPONSE          (0),
		.USE_READRESPONSE           (0),
		.USE_CLKEN                  (0),
		.AV_CONSTANT_BURST_BEHAVIOR (1),
		.AV_BURST_LINEWRAP          (0),
		.AV_BURST_BNDR_ONLY         (0),
		.AV_MAX_PENDING_READS       (4),
		.AV_MAX_PENDING_WRITES      (0),
		.AV_FIX_READ_LATENCY        (0),
		.AV_READ_WAIT_TIME          (0),
		.AV_WRITE_WAIT_TIME         (0),
		.REGISTER_WAITREQUEST       (0),
		.AV_REGISTERINCOMINGSIGNALS (0),
		.VHDL_ID                    (0)
	) fpga_mem_inst_mrx_bfm (
		.clk                      (fpga_mem_inst_afi_clk_clk),              //       clk.clk
		.reset                    (rst_controller_reset_out_reset),         // clk_reset.reset
		.avm_address              (fpga_mem_inst_mrx_bfm_m0_address),       //        m0.address
		.avm_burstcount           (fpga_mem_inst_mrx_bfm_m0_burstcount),    //          .burstcount
		.avm_readdata             (fpga_mem_inst_mrx_bfm_m0_readdata),      //          .readdata
		.avm_writedata            (fpga_mem_inst_mrx_bfm_m0_writedata),     //          .writedata
		.avm_waitrequest          (fpga_mem_inst_mrx_bfm_m0_waitrequest),   //          .waitrequest
		.avm_write                (fpga_mem_inst_mrx_bfm_m0_write),         //          .write
		.avm_read                 (fpga_mem_inst_mrx_bfm_m0_read),          //          .read
		.avm_byteenable           (fpga_mem_inst_mrx_bfm_m0_byteenable),    //          .byteenable
		.avm_readdatavalid        (fpga_mem_inst_mrx_bfm_m0_readdatavalid), //          .readdatavalid
		.avm_debugaccess          (fpga_mem_inst_mrx_bfm_m0_debugaccess),   //          .debugaccess
		.avm_begintransfer        (),                                       // (terminated)
		.avm_beginbursttransfer   (),                                       // (terminated)
		.avm_arbiterlock          (),                                       // (terminated)
		.avm_lock                 (),                                       // (terminated)
		.avm_transactionid        (),                                       // (terminated)
		.avm_readid               (8'b00000000),                            // (terminated)
		.avm_writeid              (8'b00000000),                            // (terminated)
		.avm_clken                (),                                       // (terminated)
		.avm_response             (2'b00),                                  // (terminated)
		.avm_writeresponserequest (),                                       // (terminated)
		.avm_writeresponsevalid   (1'b0),                                   // (terminated)
		.avm_readresponse         (1'b0),                                   // (terminated)
		.avm_writeresponse        (1'b0)                                    // (terminated)
	);

	altera_avalon_mm_master_bfm #(
		.AV_ADDRESS_W               (26),
		.AV_SYMBOL_W                (8),
		.AV_NUMSYMBOLS              (16),
		.AV_BURSTCOUNT_W            (6),
		.AV_READRESPONSE_W          (1),
		.AV_WRITERESPONSE_W         (1),
		.USE_READ                   (1),
		.USE_WRITE                  (1),
		.USE_ADDRESS                (1),
		.USE_BYTE_ENABLE            (1),
		.USE_BURSTCOUNT             (1),
		.USE_READ_DATA              (1),
		.USE_READ_DATA_VALID        (1),
		.USE_WRITE_DATA             (1),
		.USE_BEGIN_TRANSFER         (0),
		.USE_BEGIN_BURST_TRANSFER   (0),
		.USE_WAIT_REQUEST           (1),
		.USE_TRANSACTIONID          (0),
		.USE_WRITERESPONSE          (0),
		.USE_READRESPONSE           (0),
		.USE_CLKEN                  (0),
		.AV_CONSTANT_BURST_BEHAVIOR (1),
		.AV_BURST_LINEWRAP          (0),
		.AV_BURST_BNDR_ONLY         (0),
		.AV_MAX_PENDING_READS       (4),
		.AV_MAX_PENDING_WRITES      (0),
		.AV_FIX_READ_LATENCY        (0),
		.AV_READ_WAIT_TIME          (0),
		.AV_WRITE_WAIT_TIME         (0),
		.REGISTER_WAITREQUEST       (0),
		.AV_REGISTERINCOMINGSIGNALS (0),
		.VHDL_ID                    (1)
	) fpga_mem_inst_mr0_bfm (
		.clk                      (fpga_mem_inst_afi_clk_clk),              //       clk.clk
		.reset                    (rst_controller_reset_out_reset),         // clk_reset.reset
		.avm_address              (fpga_mem_inst_mr0_bfm_m0_address),       //        m0.address
		.avm_burstcount           (fpga_mem_inst_mr0_bfm_m0_burstcount),    //          .burstcount
		.avm_readdata             (fpga_mem_inst_mr0_bfm_m0_readdata),      //          .readdata
		.avm_writedata            (fpga_mem_inst_mr0_bfm_m0_writedata),     //          .writedata
		.avm_waitrequest          (fpga_mem_inst_mr0_bfm_m0_waitrequest),   //          .waitrequest
		.avm_write                (fpga_mem_inst_mr0_bfm_m0_write),         //          .write
		.avm_read                 (fpga_mem_inst_mr0_bfm_m0_read),          //          .read
		.avm_byteenable           (fpga_mem_inst_mr0_bfm_m0_byteenable),    //          .byteenable
		.avm_readdatavalid        (fpga_mem_inst_mr0_bfm_m0_readdatavalid), //          .readdatavalid
		.avm_debugaccess          (fpga_mem_inst_mr0_bfm_m0_debugaccess),   //          .debugaccess
		.avm_begintransfer        (),                                       // (terminated)
		.avm_beginbursttransfer   (),                                       // (terminated)
		.avm_arbiterlock          (),                                       // (terminated)
		.avm_lock                 (),                                       // (terminated)
		.avm_transactionid        (),                                       // (terminated)
		.avm_readid               (8'b00000000),                            // (terminated)
		.avm_writeid              (8'b00000000),                            // (terminated)
		.avm_clken                (),                                       // (terminated)
		.avm_response             (2'b00),                                  // (terminated)
		.avm_writeresponserequest (),                                       // (terminated)
		.avm_writeresponsevalid   (1'b0),                                   // (terminated)
		.avm_readresponse         (1'b0),                                   // (terminated)
		.avm_writeresponse        (1'b0)                                    // (terminated)
	);

	altera_avalon_mm_master_bfm #(
		.AV_ADDRESS_W               (26),
		.AV_SYMBOL_W                (8),
		.AV_NUMSYMBOLS              (16),
		.AV_BURSTCOUNT_W            (6),
		.AV_READRESPONSE_W          (1),
		.AV_WRITERESPONSE_W         (1),
		.USE_READ                   (1),
		.USE_WRITE                  (1),
		.USE_ADDRESS                (1),
		.USE_BYTE_ENABLE            (1),
		.USE_BURSTCOUNT             (1),
		.USE_READ_DATA              (1),
		.USE_READ_DATA_VALID        (1),
		.USE_WRITE_DATA             (1),
		.USE_BEGIN_TRANSFER         (0),
		.USE_BEGIN_BURST_TRANSFER   (0),
		.USE_WAIT_REQUEST           (1),
		.USE_TRANSACTIONID          (0),
		.USE_WRITERESPONSE          (0),
		.USE_READRESPONSE           (0),
		.USE_CLKEN                  (0),
		.AV_CONSTANT_BURST_BEHAVIOR (1),
		.AV_BURST_LINEWRAP          (0),
		.AV_BURST_BNDR_ONLY         (0),
		.AV_MAX_PENDING_READS       (4),
		.AV_MAX_PENDING_WRITES      (0),
		.AV_FIX_READ_LATENCY        (0),
		.AV_READ_WAIT_TIME          (0),
		.AV_WRITE_WAIT_TIME         (0),
		.REGISTER_WAITREQUEST       (0),
		.AV_REGISTERINCOMINGSIGNALS (0),
		.VHDL_ID                    (2)
	) fpga_mem_inst_mr1_bfm (
		.clk                      (fpga_mem_inst_afi_clk_clk),              //       clk.clk
		.reset                    (rst_controller_reset_out_reset),         // clk_reset.reset
		.avm_address              (fpga_mem_inst_mr1_bfm_m0_address),       //        m0.address
		.avm_burstcount           (fpga_mem_inst_mr1_bfm_m0_burstcount),    //          .burstcount
		.avm_readdata             (fpga_mem_inst_mr1_bfm_m0_readdata),      //          .readdata
		.avm_writedata            (fpga_mem_inst_mr1_bfm_m0_writedata),     //          .writedata
		.avm_waitrequest          (fpga_mem_inst_mr1_bfm_m0_waitrequest),   //          .waitrequest
		.avm_write                (fpga_mem_inst_mr1_bfm_m0_write),         //          .write
		.avm_read                 (fpga_mem_inst_mr1_bfm_m0_read),          //          .read
		.avm_byteenable           (fpga_mem_inst_mr1_bfm_m0_byteenable),    //          .byteenable
		.avm_readdatavalid        (fpga_mem_inst_mr1_bfm_m0_readdatavalid), //          .readdatavalid
		.avm_debugaccess          (fpga_mem_inst_mr1_bfm_m0_debugaccess),   //          .debugaccess
		.avm_begintransfer        (),                                       // (terminated)
		.avm_beginbursttransfer   (),                                       // (terminated)
		.avm_arbiterlock          (),                                       // (terminated)
		.avm_lock                 (),                                       // (terminated)
		.avm_transactionid        (),                                       // (terminated)
		.avm_readid               (8'b00000000),                            // (terminated)
		.avm_writeid              (8'b00000000),                            // (terminated)
		.avm_clken                (),                                       // (terminated)
		.avm_response             (2'b00),                                  // (terminated)
		.avm_writeresponserequest (),                                       // (terminated)
		.avm_writeresponsevalid   (1'b0),                                   // (terminated)
		.avm_readresponse         (1'b0),                                   // (terminated)
		.avm_writeresponse        (1'b0)                                    // (terminated)
	);

	altera_avalon_mm_master_bfm #(
		.AV_ADDRESS_W               (26),
		.AV_SYMBOL_W                (8),
		.AV_NUMSYMBOLS              (16),
		.AV_BURSTCOUNT_W            (6),
		.AV_READRESPONSE_W          (1),
		.AV_WRITERESPONSE_W         (1),
		.USE_READ                   (1),
		.USE_WRITE                  (1),
		.USE_ADDRESS                (1),
		.USE_BYTE_ENABLE            (1),
		.USE_BURSTCOUNT             (1),
		.USE_READ_DATA              (1),
		.USE_READ_DATA_VALID        (1),
		.USE_WRITE_DATA             (1),
		.USE_BEGIN_TRANSFER         (0),
		.USE_BEGIN_BURST_TRANSFER   (0),
		.USE_WAIT_REQUEST           (1),
		.USE_TRANSACTIONID          (0),
		.USE_WRITERESPONSE          (0),
		.USE_READRESPONSE           (0),
		.USE_CLKEN                  (0),
		.AV_CONSTANT_BURST_BEHAVIOR (1),
		.AV_BURST_LINEWRAP          (0),
		.AV_BURST_BNDR_ONLY         (0),
		.AV_MAX_PENDING_READS       (4),
		.AV_MAX_PENDING_WRITES      (0),
		.AV_FIX_READ_LATENCY        (0),
		.AV_READ_WAIT_TIME          (0),
		.AV_WRITE_WAIT_TIME         (0),
		.REGISTER_WAITREQUEST       (0),
		.AV_REGISTERINCOMINGSIGNALS (0),
		.VHDL_ID                    (3)
	) fpga_mem_inst_mr2_bfm (
		.clk                      (fpga_mem_inst_afi_clk_clk),              //       clk.clk
		.reset                    (rst_controller_reset_out_reset),         // clk_reset.reset
		.avm_address              (fpga_mem_inst_mr2_bfm_m0_address),       //        m0.address
		.avm_burstcount           (fpga_mem_inst_mr2_bfm_m0_burstcount),    //          .burstcount
		.avm_readdata             (fpga_mem_inst_mr2_bfm_m0_readdata),      //          .readdata
		.avm_writedata            (fpga_mem_inst_mr2_bfm_m0_writedata),     //          .writedata
		.avm_waitrequest          (fpga_mem_inst_mr2_bfm_m0_waitrequest),   //          .waitrequest
		.avm_write                (fpga_mem_inst_mr2_bfm_m0_write),         //          .write
		.avm_read                 (fpga_mem_inst_mr2_bfm_m0_read),          //          .read
		.avm_byteenable           (fpga_mem_inst_mr2_bfm_m0_byteenable),    //          .byteenable
		.avm_readdatavalid        (fpga_mem_inst_mr2_bfm_m0_readdatavalid), //          .readdatavalid
		.avm_debugaccess          (fpga_mem_inst_mr2_bfm_m0_debugaccess),   //          .debugaccess
		.avm_begintransfer        (),                                       // (terminated)
		.avm_beginbursttransfer   (),                                       // (terminated)
		.avm_arbiterlock          (),                                       // (terminated)
		.avm_lock                 (),                                       // (terminated)
		.avm_transactionid        (),                                       // (terminated)
		.avm_readid               (8'b00000000),                            // (terminated)
		.avm_writeid              (8'b00000000),                            // (terminated)
		.avm_clken                (),                                       // (terminated)
		.avm_response             (2'b00),                                  // (terminated)
		.avm_writeresponserequest (),                                       // (terminated)
		.avm_writeresponsevalid   (1'b0),                                   // (terminated)
		.avm_readresponse         (1'b0),                                   // (terminated)
		.avm_writeresponse        (1'b0)                                    // (terminated)
	);

	altera_avalon_mm_master_bfm #(
		.AV_ADDRESS_W               (26),
		.AV_SYMBOL_W                (8),
		.AV_NUMSYMBOLS              (16),
		.AV_BURSTCOUNT_W            (6),
		.AV_READRESPONSE_W          (1),
		.AV_WRITERESPONSE_W         (1),
		.USE_READ                   (1),
		.USE_WRITE                  (1),
		.USE_ADDRESS                (1),
		.USE_BYTE_ENABLE            (1),
		.USE_BURSTCOUNT             (1),
		.USE_READ_DATA              (1),
		.USE_READ_DATA_VALID        (1),
		.USE_WRITE_DATA             (1),
		.USE_BEGIN_TRANSFER         (0),
		.USE_BEGIN_BURST_TRANSFER   (0),
		.USE_WAIT_REQUEST           (1),
		.USE_TRANSACTIONID          (0),
		.USE_WRITERESPONSE          (0),
		.USE_READRESPONSE           (0),
		.USE_CLKEN                  (0),
		.AV_CONSTANT_BURST_BEHAVIOR (1),
		.AV_BURST_LINEWRAP          (0),
		.AV_BURST_BNDR_ONLY         (0),
		.AV_MAX_PENDING_READS       (4),
		.AV_MAX_PENDING_WRITES      (0),
		.AV_FIX_READ_LATENCY        (0),
		.AV_READ_WAIT_TIME          (0),
		.AV_WRITE_WAIT_TIME         (0),
		.REGISTER_WAITREQUEST       (0),
		.AV_REGISTERINCOMINGSIGNALS (0),
		.VHDL_ID                    (4)
	) fpga_mem_inst_mr3_bfm (
		.clk                      (fpga_mem_inst_afi_clk_clk),              //       clk.clk
		.reset                    (rst_controller_reset_out_reset),         // clk_reset.reset
		.avm_address              (fpga_mem_inst_mr3_bfm_m0_address),       //        m0.address
		.avm_burstcount           (fpga_mem_inst_mr3_bfm_m0_burstcount),    //          .burstcount
		.avm_readdata             (fpga_mem_inst_mr3_bfm_m0_readdata),      //          .readdata
		.avm_writedata            (fpga_mem_inst_mr3_bfm_m0_writedata),     //          .writedata
		.avm_waitrequest          (fpga_mem_inst_mr3_bfm_m0_waitrequest),   //          .waitrequest
		.avm_write                (fpga_mem_inst_mr3_bfm_m0_write),         //          .write
		.avm_read                 (fpga_mem_inst_mr3_bfm_m0_read),          //          .read
		.avm_byteenable           (fpga_mem_inst_mr3_bfm_m0_byteenable),    //          .byteenable
		.avm_readdatavalid        (fpga_mem_inst_mr3_bfm_m0_readdatavalid), //          .readdatavalid
		.avm_debugaccess          (fpga_mem_inst_mr3_bfm_m0_debugaccess),   //          .debugaccess
		.avm_begintransfer        (),                                       // (terminated)
		.avm_beginbursttransfer   (),                                       // (terminated)
		.avm_arbiterlock          (),                                       // (terminated)
		.avm_lock                 (),                                       // (terminated)
		.avm_transactionid        (),                                       // (terminated)
		.avm_readid               (8'b00000000),                            // (terminated)
		.avm_writeid              (8'b00000000),                            // (terminated)
		.avm_clken                (),                                       // (terminated)
		.avm_response             (2'b00),                                  // (terminated)
		.avm_writeresponserequest (),                                       // (terminated)
		.avm_writeresponsevalid   (1'b0),                                   // (terminated)
		.avm_readresponse         (1'b0),                                   // (terminated)
		.avm_writeresponse        (1'b0)                                    // (terminated)
	);

	altera_avalon_mm_master_bfm #(
		.AV_ADDRESS_W               (26),
		.AV_SYMBOL_W                (8),
		.AV_NUMSYMBOLS              (16),
		.AV_BURSTCOUNT_W            (6),
		.AV_READRESPONSE_W          (1),
		.AV_WRITERESPONSE_W         (1),
		.USE_READ                   (1),
		.USE_WRITE                  (1),
		.USE_ADDRESS                (1),
		.USE_BYTE_ENABLE            (1),
		.USE_BURSTCOUNT             (1),
		.USE_READ_DATA              (1),
		.USE_READ_DATA_VALID        (1),
		.USE_WRITE_DATA             (1),
		.USE_BEGIN_TRANSFER         (0),
		.USE_BEGIN_BURST_TRANSFER   (0),
		.USE_WAIT_REQUEST           (1),
		.USE_TRANSACTIONID          (0),
		.USE_WRITERESPONSE          (0),
		.USE_READRESPONSE           (0),
		.USE_CLKEN                  (0),
		.AV_CONSTANT_BURST_BEHAVIOR (1),
		.AV_BURST_LINEWRAP          (0),
		.AV_BURST_BNDR_ONLY         (0),
		.AV_MAX_PENDING_READS       (4),
		.AV_MAX_PENDING_WRITES      (0),
		.AV_FIX_READ_LATENCY        (0),
		.AV_READ_WAIT_TIME          (0),
		.AV_WRITE_WAIT_TIME         (0),
		.REGISTER_WAITREQUEST       (0),
		.AV_REGISTERINCOMINGSIGNALS (0),
		.VHDL_ID                    (5)
	) fpga_mem_inst_mwx_bfm (
		.clk                      (fpga_mem_inst_afi_clk_clk),              //       clk.clk
		.reset                    (rst_controller_reset_out_reset),         // clk_reset.reset
		.avm_address              (fpga_mem_inst_mwx_bfm_m0_address),       //        m0.address
		.avm_burstcount           (fpga_mem_inst_mwx_bfm_m0_burstcount),    //          .burstcount
		.avm_readdata             (fpga_mem_inst_mwx_bfm_m0_readdata),      //          .readdata
		.avm_writedata            (fpga_mem_inst_mwx_bfm_m0_writedata),     //          .writedata
		.avm_waitrequest          (fpga_mem_inst_mwx_bfm_m0_waitrequest),   //          .waitrequest
		.avm_write                (fpga_mem_inst_mwx_bfm_m0_write),         //          .write
		.avm_read                 (fpga_mem_inst_mwx_bfm_m0_read),          //          .read
		.avm_byteenable           (fpga_mem_inst_mwx_bfm_m0_byteenable),    //          .byteenable
		.avm_readdatavalid        (fpga_mem_inst_mwx_bfm_m0_readdatavalid), //          .readdatavalid
		.avm_debugaccess          (fpga_mem_inst_mwx_bfm_m0_debugaccess),   //          .debugaccess
		.avm_begintransfer        (),                                       // (terminated)
		.avm_beginbursttransfer   (),                                       // (terminated)
		.avm_arbiterlock          (),                                       // (terminated)
		.avm_lock                 (),                                       // (terminated)
		.avm_transactionid        (),                                       // (terminated)
		.avm_readid               (8'b00000000),                            // (terminated)
		.avm_writeid              (8'b00000000),                            // (terminated)
		.avm_clken                (),                                       // (terminated)
		.avm_response             (2'b00),                                  // (terminated)
		.avm_writeresponserequest (),                                       // (terminated)
		.avm_writeresponsevalid   (1'b0),                                   // (terminated)
		.avm_readresponse         (1'b0),                                   // (terminated)
		.avm_writeresponse        (1'b0)                                    // (terminated)
	);

	altera_avalon_mm_master_bfm #(
		.AV_ADDRESS_W               (26),
		.AV_SYMBOL_W                (8),
		.AV_NUMSYMBOLS              (16),
		.AV_BURSTCOUNT_W            (6),
		.AV_READRESPONSE_W          (1),
		.AV_WRITERESPONSE_W         (1),
		.USE_READ                   (1),
		.USE_WRITE                  (1),
		.USE_ADDRESS                (1),
		.USE_BYTE_ENABLE            (1),
		.USE_BURSTCOUNT             (1),
		.USE_READ_DATA              (1),
		.USE_READ_DATA_VALID        (1),
		.USE_WRITE_DATA             (1),
		.USE_BEGIN_TRANSFER         (0),
		.USE_BEGIN_BURST_TRANSFER   (0),
		.USE_WAIT_REQUEST           (1),
		.USE_TRANSACTIONID          (0),
		.USE_WRITERESPONSE          (0),
		.USE_READRESPONSE           (0),
		.USE_CLKEN                  (0),
		.AV_CONSTANT_BURST_BEHAVIOR (1),
		.AV_BURST_LINEWRAP          (0),
		.AV_BURST_BNDR_ONLY         (0),
		.AV_MAX_PENDING_READS       (4),
		.AV_MAX_PENDING_WRITES      (0),
		.AV_FIX_READ_LATENCY        (0),
		.AV_READ_WAIT_TIME          (0),
		.AV_WRITE_WAIT_TIME         (0),
		.REGISTER_WAITREQUEST       (0),
		.AV_REGISTERINCOMINGSIGNALS (0),
		.VHDL_ID                    (6)
	) fpga_mem_inst_mw0_bfm (
		.clk                      (fpga_mem_inst_afi_clk_clk),              //       clk.clk
		.reset                    (rst_controller_reset_out_reset),         // clk_reset.reset
		.avm_address              (fpga_mem_inst_mw0_bfm_m0_address),       //        m0.address
		.avm_burstcount           (fpga_mem_inst_mw0_bfm_m0_burstcount),    //          .burstcount
		.avm_readdata             (fpga_mem_inst_mw0_bfm_m0_readdata),      //          .readdata
		.avm_writedata            (fpga_mem_inst_mw0_bfm_m0_writedata),     //          .writedata
		.avm_waitrequest          (fpga_mem_inst_mw0_bfm_m0_waitrequest),   //          .waitrequest
		.avm_write                (fpga_mem_inst_mw0_bfm_m0_write),         //          .write
		.avm_read                 (fpga_mem_inst_mw0_bfm_m0_read),          //          .read
		.avm_byteenable           (fpga_mem_inst_mw0_bfm_m0_byteenable),    //          .byteenable
		.avm_readdatavalid        (fpga_mem_inst_mw0_bfm_m0_readdatavalid), //          .readdatavalid
		.avm_debugaccess          (fpga_mem_inst_mw0_bfm_m0_debugaccess),   //          .debugaccess
		.avm_begintransfer        (),                                       // (terminated)
		.avm_beginbursttransfer   (),                                       // (terminated)
		.avm_arbiterlock          (),                                       // (terminated)
		.avm_lock                 (),                                       // (terminated)
		.avm_transactionid        (),                                       // (terminated)
		.avm_readid               (8'b00000000),                            // (terminated)
		.avm_writeid              (8'b00000000),                            // (terminated)
		.avm_clken                (),                                       // (terminated)
		.avm_response             (2'b00),                                  // (terminated)
		.avm_writeresponserequest (),                                       // (terminated)
		.avm_writeresponsevalid   (1'b0),                                   // (terminated)
		.avm_readresponse         (1'b0),                                   // (terminated)
		.avm_writeresponse        (1'b0)                                    // (terminated)
	);

	altera_avalon_mm_master_bfm #(
		.AV_ADDRESS_W               (26),
		.AV_SYMBOL_W                (8),
		.AV_NUMSYMBOLS              (16),
		.AV_BURSTCOUNT_W            (6),
		.AV_READRESPONSE_W          (1),
		.AV_WRITERESPONSE_W         (1),
		.USE_READ                   (1),
		.USE_WRITE                  (1),
		.USE_ADDRESS                (1),
		.USE_BYTE_ENABLE            (1),
		.USE_BURSTCOUNT             (1),
		.USE_READ_DATA              (1),
		.USE_READ_DATA_VALID        (1),
		.USE_WRITE_DATA             (1),
		.USE_BEGIN_TRANSFER         (0),
		.USE_BEGIN_BURST_TRANSFER   (0),
		.USE_WAIT_REQUEST           (1),
		.USE_TRANSACTIONID          (0),
		.USE_WRITERESPONSE          (0),
		.USE_READRESPONSE           (0),
		.USE_CLKEN                  (0),
		.AV_CONSTANT_BURST_BEHAVIOR (1),
		.AV_BURST_LINEWRAP          (0),
		.AV_BURST_BNDR_ONLY         (0),
		.AV_MAX_PENDING_READS       (4),
		.AV_MAX_PENDING_WRITES      (0),
		.AV_FIX_READ_LATENCY        (0),
		.AV_READ_WAIT_TIME          (0),
		.AV_WRITE_WAIT_TIME         (0),
		.REGISTER_WAITREQUEST       (0),
		.AV_REGISTERINCOMINGSIGNALS (0),
		.VHDL_ID                    (7)
	) fpga_mem_inst_mw1_bfm (
		.clk                      (fpga_mem_inst_afi_clk_clk),              //       clk.clk
		.reset                    (rst_controller_reset_out_reset),         // clk_reset.reset
		.avm_address              (fpga_mem_inst_mw1_bfm_m0_address),       //        m0.address
		.avm_burstcount           (fpga_mem_inst_mw1_bfm_m0_burstcount),    //          .burstcount
		.avm_readdata             (fpga_mem_inst_mw1_bfm_m0_readdata),      //          .readdata
		.avm_writedata            (fpga_mem_inst_mw1_bfm_m0_writedata),     //          .writedata
		.avm_waitrequest          (fpga_mem_inst_mw1_bfm_m0_waitrequest),   //          .waitrequest
		.avm_write                (fpga_mem_inst_mw1_bfm_m0_write),         //          .write
		.avm_read                 (fpga_mem_inst_mw1_bfm_m0_read),          //          .read
		.avm_byteenable           (fpga_mem_inst_mw1_bfm_m0_byteenable),    //          .byteenable
		.avm_readdatavalid        (fpga_mem_inst_mw1_bfm_m0_readdatavalid), //          .readdatavalid
		.avm_debugaccess          (fpga_mem_inst_mw1_bfm_m0_debugaccess),   //          .debugaccess
		.avm_begintransfer        (),                                       // (terminated)
		.avm_beginbursttransfer   (),                                       // (terminated)
		.avm_arbiterlock          (),                                       // (terminated)
		.avm_lock                 (),                                       // (terminated)
		.avm_transactionid        (),                                       // (terminated)
		.avm_readid               (8'b00000000),                            // (terminated)
		.avm_writeid              (8'b00000000),                            // (terminated)
		.avm_clken                (),                                       // (terminated)
		.avm_response             (2'b00),                                  // (terminated)
		.avm_writeresponserequest (),                                       // (terminated)
		.avm_writeresponsevalid   (1'b0),                                   // (terminated)
		.avm_readresponse         (1'b0),                                   // (terminated)
		.avm_writeresponse        (1'b0)                                    // (terminated)
	);

	altera_avalon_mm_master_bfm #(
		.AV_ADDRESS_W               (26),
		.AV_SYMBOL_W                (8),
		.AV_NUMSYMBOLS              (16),
		.AV_BURSTCOUNT_W            (6),
		.AV_READRESPONSE_W          (1),
		.AV_WRITERESPONSE_W         (1),
		.USE_READ                   (1),
		.USE_WRITE                  (1),
		.USE_ADDRESS                (1),
		.USE_BYTE_ENABLE            (1),
		.USE_BURSTCOUNT             (1),
		.USE_READ_DATA              (1),
		.USE_READ_DATA_VALID        (1),
		.USE_WRITE_DATA             (1),
		.USE_BEGIN_TRANSFER         (0),
		.USE_BEGIN_BURST_TRANSFER   (0),
		.USE_WAIT_REQUEST           (1),
		.USE_TRANSACTIONID          (0),
		.USE_WRITERESPONSE          (0),
		.USE_READRESPONSE           (0),
		.USE_CLKEN                  (0),
		.AV_CONSTANT_BURST_BEHAVIOR (1),
		.AV_BURST_LINEWRAP          (0),
		.AV_BURST_BNDR_ONLY         (0),
		.AV_MAX_PENDING_READS       (4),
		.AV_MAX_PENDING_WRITES      (0),
		.AV_FIX_READ_LATENCY        (0),
		.AV_READ_WAIT_TIME          (0),
		.AV_WRITE_WAIT_TIME         (0),
		.REGISTER_WAITREQUEST       (0),
		.AV_REGISTERINCOMINGSIGNALS (0),
		.VHDL_ID                    (8)
	) fpga_mem_inst_mw2_bfm (
		.clk                      (fpga_mem_inst_afi_clk_clk),              //       clk.clk
		.reset                    (rst_controller_reset_out_reset),         // clk_reset.reset
		.avm_address              (fpga_mem_inst_mw2_bfm_m0_address),       //        m0.address
		.avm_burstcount           (fpga_mem_inst_mw2_bfm_m0_burstcount),    //          .burstcount
		.avm_readdata             (fpga_mem_inst_mw2_bfm_m0_readdata),      //          .readdata
		.avm_writedata            (fpga_mem_inst_mw2_bfm_m0_writedata),     //          .writedata
		.avm_waitrequest          (fpga_mem_inst_mw2_bfm_m0_waitrequest),   //          .waitrequest
		.avm_write                (fpga_mem_inst_mw2_bfm_m0_write),         //          .write
		.avm_read                 (fpga_mem_inst_mw2_bfm_m0_read),          //          .read
		.avm_byteenable           (fpga_mem_inst_mw2_bfm_m0_byteenable),    //          .byteenable
		.avm_readdatavalid        (fpga_mem_inst_mw2_bfm_m0_readdatavalid), //          .readdatavalid
		.avm_debugaccess          (fpga_mem_inst_mw2_bfm_m0_debugaccess),   //          .debugaccess
		.avm_begintransfer        (),                                       // (terminated)
		.avm_beginbursttransfer   (),                                       // (terminated)
		.avm_arbiterlock          (),                                       // (terminated)
		.avm_lock                 (),                                       // (terminated)
		.avm_transactionid        (),                                       // (terminated)
		.avm_readid               (8'b00000000),                            // (terminated)
		.avm_writeid              (8'b00000000),                            // (terminated)
		.avm_clken                (),                                       // (terminated)
		.avm_response             (2'b00),                                  // (terminated)
		.avm_writeresponserequest (),                                       // (terminated)
		.avm_writeresponsevalid   (1'b0),                                   // (terminated)
		.avm_readresponse         (1'b0),                                   // (terminated)
		.avm_writeresponse        (1'b0)                                    // (terminated)
	);

	altera_avalon_mm_master_bfm #(
		.AV_ADDRESS_W               (26),
		.AV_SYMBOL_W                (8),
		.AV_NUMSYMBOLS              (16),
		.AV_BURSTCOUNT_W            (6),
		.AV_READRESPONSE_W          (1),
		.AV_WRITERESPONSE_W         (1),
		.USE_READ                   (1),
		.USE_WRITE                  (1),
		.USE_ADDRESS                (1),
		.USE_BYTE_ENABLE            (1),
		.USE_BURSTCOUNT             (1),
		.USE_READ_DATA              (1),
		.USE_READ_DATA_VALID        (1),
		.USE_WRITE_DATA             (1),
		.USE_BEGIN_TRANSFER         (0),
		.USE_BEGIN_BURST_TRANSFER   (0),
		.USE_WAIT_REQUEST           (1),
		.USE_TRANSACTIONID          (0),
		.USE_WRITERESPONSE          (0),
		.USE_READRESPONSE           (0),
		.USE_CLKEN                  (0),
		.AV_CONSTANT_BURST_BEHAVIOR (1),
		.AV_BURST_LINEWRAP          (0),
		.AV_BURST_BNDR_ONLY         (0),
		.AV_MAX_PENDING_READS       (4),
		.AV_MAX_PENDING_WRITES      (0),
		.AV_FIX_READ_LATENCY        (0),
		.AV_READ_WAIT_TIME          (0),
		.AV_WRITE_WAIT_TIME         (0),
		.REGISTER_WAITREQUEST       (0),
		.AV_REGISTERINCOMINGSIGNALS (0),
		.VHDL_ID                    (9)
	) fpga_mem_inst_mw3_bfm (
		.clk                      (fpga_mem_inst_afi_clk_clk),              //       clk.clk
		.reset                    (rst_controller_reset_out_reset),         // clk_reset.reset
		.avm_address              (fpga_mem_inst_mw3_bfm_m0_address),       //        m0.address
		.avm_burstcount           (fpga_mem_inst_mw3_bfm_m0_burstcount),    //          .burstcount
		.avm_readdata             (fpga_mem_inst_mw3_bfm_m0_readdata),      //          .readdata
		.avm_writedata            (fpga_mem_inst_mw3_bfm_m0_writedata),     //          .writedata
		.avm_waitrequest          (fpga_mem_inst_mw3_bfm_m0_waitrequest),   //          .waitrequest
		.avm_write                (fpga_mem_inst_mw3_bfm_m0_write),         //          .write
		.avm_read                 (fpga_mem_inst_mw3_bfm_m0_read),          //          .read
		.avm_byteenable           (fpga_mem_inst_mw3_bfm_m0_byteenable),    //          .byteenable
		.avm_readdatavalid        (fpga_mem_inst_mw3_bfm_m0_readdatavalid), //          .readdatavalid
		.avm_debugaccess          (fpga_mem_inst_mw3_bfm_m0_debugaccess),   //          .debugaccess
		.avm_begintransfer        (),                                       // (terminated)
		.avm_beginbursttransfer   (),                                       // (terminated)
		.avm_arbiterlock          (),                                       // (terminated)
		.avm_lock                 (),                                       // (terminated)
		.avm_transactionid        (),                                       // (terminated)
		.avm_readid               (8'b00000000),                            // (terminated)
		.avm_writeid              (8'b00000000),                            // (terminated)
		.avm_clken                (),                                       // (terminated)
		.avm_response             (2'b00),                                  // (terminated)
		.avm_writeresponserequest (),                                       // (terminated)
		.avm_writeresponsevalid   (1'b0),                                   // (terminated)
		.avm_readresponse         (1'b0),                                   // (terminated)
		.avm_writeresponse        (1'b0)                                    // (terminated)
	);

	altera_avalon_mm_master_bfm #(
		.AV_ADDRESS_W               (26),
		.AV_SYMBOL_W                (8),
		.AV_NUMSYMBOLS              (16),
		.AV_BURSTCOUNT_W            (6),
		.AV_READRESPONSE_W          (1),
		.AV_WRITERESPONSE_W         (1),
		.USE_READ                   (1),
		.USE_WRITE                  (1),
		.USE_ADDRESS                (1),
		.USE_BYTE_ENABLE            (1),
		.USE_BURSTCOUNT             (1),
		.USE_READ_DATA              (1),
		.USE_READ_DATA_VALID        (1),
		.USE_WRITE_DATA             (1),
		.USE_BEGIN_TRANSFER         (0),
		.USE_BEGIN_BURST_TRANSFER   (0),
		.USE_WAIT_REQUEST           (1),
		.USE_TRANSACTIONID          (0),
		.USE_WRITERESPONSE          (0),
		.USE_READRESPONSE           (0),
		.USE_CLKEN                  (0),
		.AV_CONSTANT_BURST_BEHAVIOR (1),
		.AV_BURST_LINEWRAP          (0),
		.AV_BURST_BNDR_ONLY         (0),
		.AV_MAX_PENDING_READS       (4),
		.AV_MAX_PENDING_WRITES      (0),
		.AV_FIX_READ_LATENCY        (0),
		.AV_READ_WAIT_TIME          (0),
		.AV_WRITE_WAIT_TIME         (0),
		.REGISTER_WAITREQUEST       (0),
		.AV_REGISTERINCOMINGSIGNALS (0),
		.VHDL_ID                    (10)
	) fpga_mem_inst_hps_bfm (
		.clk                      (fpga_mem_inst_afi_clk_clk),              //       clk.clk
		.reset                    (rst_controller_reset_out_reset),         // clk_reset.reset
		.avm_address              (fpga_mem_inst_hps_bfm_m0_address),       //        m0.address
		.avm_burstcount           (fpga_mem_inst_hps_bfm_m0_burstcount),    //          .burstcount
		.avm_readdata             (fpga_mem_inst_hps_bfm_m0_readdata),      //          .readdata
		.avm_writedata            (fpga_mem_inst_hps_bfm_m0_writedata),     //          .writedata
		.avm_waitrequest          (fpga_mem_inst_hps_bfm_m0_waitrequest),   //          .waitrequest
		.avm_write                (fpga_mem_inst_hps_bfm_m0_write),         //          .write
		.avm_read                 (fpga_mem_inst_hps_bfm_m0_read),          //          .read
		.avm_byteenable           (fpga_mem_inst_hps_bfm_m0_byteenable),    //          .byteenable
		.avm_readdatavalid        (fpga_mem_inst_hps_bfm_m0_readdatavalid), //          .readdatavalid
		.avm_debugaccess          (fpga_mem_inst_hps_bfm_m0_debugaccess),   //          .debugaccess
		.avm_begintransfer        (),                                       // (terminated)
		.avm_beginbursttransfer   (),                                       // (terminated)
		.avm_arbiterlock          (),                                       // (terminated)
		.avm_lock                 (),                                       // (terminated)
		.avm_transactionid        (),                                       // (terminated)
		.avm_readid               (8'b00000000),                            // (terminated)
		.avm_writeid              (8'b00000000),                            // (terminated)
		.avm_clken                (),                                       // (terminated)
		.avm_response             (2'b00),                                  // (terminated)
		.avm_writeresponserequest (),                                       // (terminated)
		.avm_writeresponsevalid   (1'b0),                                   // (terminated)
		.avm_readresponse         (1'b0),                                   // (terminated)
		.avm_writeresponse        (1'b0)                                    // (terminated)
	);

	alt_mem_if_ddr3_mem_model_top_ddr3_mem_if_dm_pins_en_mem_if_dqsn_en #(
		.MEM_IF_ADDR_WIDTH              (15),
		.MEM_IF_ROW_ADDR_WIDTH          (15),
		.MEM_IF_COL_ADDR_WIDTH          (10),
		.MEM_IF_CONTROL_WIDTH           (1),
		.MEM_IF_DQS_WIDTH               (4),
		.MEM_IF_CS_WIDTH                (1),
		.MEM_IF_BANKADDR_WIDTH          (3),
		.MEM_IF_DQ_WIDTH                (32),
		.MEM_IF_CK_WIDTH                (1),
		.MEM_IF_CLK_EN_WIDTH            (1),
		.DEVICE_WIDTH                   (1),
		.MEM_TRCD                       (5),
		.MEM_TRTP                       (4),
		.MEM_DQS_TO_CLK_CAPTURE_DELAY   (450),
		.MEM_CLK_TO_DQS_CAPTURE_DELAY   (100000),
		.MEM_IF_ODT_WIDTH               (1),
		.MEM_MIRROR_ADDRESSING_DEC      (0),
		.MEM_REGDIMM_ENABLED            (0),
		.MEM_LRDIMM_ENABLED             (0),
		.DEVICE_DEPTH                   (1),
		.MEM_NUMBER_OF_DIMMS            (1),
		.MEM_NUMBER_OF_RANKS_PER_DIMM   (1),
		.MEM_RANK_MULTIPLICATION_FACTOR (1),
		.MEM_GUARANTEED_WRITE_INIT      (0),
		.MEM_VERBOSE                    (1),
		.REFRESH_BURST_VALIDATION       (0),
		.MEM_INIT_EN                    (0),
		.MEM_INIT_FILE                  (""),
		.DAT_DATA_WIDTH                 (32)
	) mem_if_ddr3_emif_0_mem_model (
		.mem_a       (fpga_mem_inst_memory_0_mem_a),       // memory.mem_a
		.mem_ba      (fpga_mem_inst_memory_0_mem_ba),      //       .mem_ba
		.mem_ck      (fpga_mem_inst_memory_0_mem_ck),      //       .mem_ck
		.mem_ck_n    (fpga_mem_inst_memory_0_mem_ck_n),    //       .mem_ck_n
		.mem_cke     (fpga_mem_inst_memory_0_mem_cke),     //       .mem_cke
		.mem_cs_n    (fpga_mem_inst_memory_0_mem_cs_n),    //       .mem_cs_n
		.mem_dm      (fpga_mem_inst_memory_0_mem_dm),      //       .mem_dm
		.mem_ras_n   (fpga_mem_inst_memory_0_mem_ras_n),   //       .mem_ras_n
		.mem_cas_n   (fpga_mem_inst_memory_0_mem_cas_n),   //       .mem_cas_n
		.mem_we_n    (fpga_mem_inst_memory_0_mem_we_n),    //       .mem_we_n
		.mem_reset_n (fpga_mem_inst_memory_0_mem_reset_n), //       .mem_reset_n
		.mem_dq      (fpga_mem_inst_memory_0_mem_dq),      //       .mem_dq
		.mem_dqs     (fpga_mem_inst_memory_0_mem_dqs),     //       .mem_dqs
		.mem_dqs_n   (fpga_mem_inst_memory_0_mem_dqs_n),   //       .mem_dqs_n
		.mem_odt     (fpga_mem_inst_memory_0_mem_odt)      //       .mem_odt
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~fpga_mem_inst_reset_bfm_reset_reset), // reset_in0.reset
		.clk            (fpga_mem_inst_afi_clk_clk),            //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),       // reset_out.reset
		.reset_req      (),                                     // (terminated)
		.reset_req_in0  (1'b0),                                 // (terminated)
		.reset_in1      (1'b0),                                 // (terminated)
		.reset_req_in1  (1'b0),                                 // (terminated)
		.reset_in2      (1'b0),                                 // (terminated)
		.reset_req_in2  (1'b0),                                 // (terminated)
		.reset_in3      (1'b0),                                 // (terminated)
		.reset_req_in3  (1'b0),                                 // (terminated)
		.reset_in4      (1'b0),                                 // (terminated)
		.reset_req_in4  (1'b0),                                 // (terminated)
		.reset_in5      (1'b0),                                 // (terminated)
		.reset_req_in5  (1'b0),                                 // (terminated)
		.reset_in6      (1'b0),                                 // (terminated)
		.reset_req_in6  (1'b0),                                 // (terminated)
		.reset_in7      (1'b0),                                 // (terminated)
		.reset_req_in7  (1'b0),                                 // (terminated)
		.reset_in8      (1'b0),                                 // (terminated)
		.reset_req_in8  (1'b0),                                 // (terminated)
		.reset_in9      (1'b0),                                 // (terminated)
		.reset_req_in9  (1'b0),                                 // (terminated)
		.reset_in10     (1'b0),                                 // (terminated)
		.reset_req_in10 (1'b0),                                 // (terminated)
		.reset_in11     (1'b0),                                 // (terminated)
		.reset_req_in11 (1'b0),                                 // (terminated)
		.reset_in12     (1'b0),                                 // (terminated)
		.reset_req_in12 (1'b0),                                 // (terminated)
		.reset_in13     (1'b0),                                 // (terminated)
		.reset_req_in13 (1'b0),                                 // (terminated)
		.reset_in14     (1'b0),                                 // (terminated)
		.reset_req_in14 (1'b0),                                 // (terminated)
		.reset_in15     (1'b0),                                 // (terminated)
		.reset_req_in15 (1'b0)                                  // (terminated)
	);

endmodule
