// fpga_mem.v

// Generated using ACDS version 13.1 162 at 2015.07.03.12:59:18

`timescale 1 ps / 1 ps
module fpga_mem (
		input  wire         clk_clk,                                                  //                            clk.clk
		input  wire         reset_reset_n,                                            //                          reset.reset_n
		output wire [14:0]  memory_0_mem_a,                                           //                       memory_0.mem_a
		output wire [2:0]   memory_0_mem_ba,                                          //                               .mem_ba
		output wire [0:0]   memory_0_mem_ck,                                          //                               .mem_ck
		output wire [0:0]   memory_0_mem_ck_n,                                        //                               .mem_ck_n
		output wire [0:0]   memory_0_mem_cke,                                         //                               .mem_cke
		output wire [0:0]   memory_0_mem_cs_n,                                        //                               .mem_cs_n
		output wire [3:0]   memory_0_mem_dm,                                          //                               .mem_dm
		output wire [0:0]   memory_0_mem_ras_n,                                       //                               .mem_ras_n
		output wire [0:0]   memory_0_mem_cas_n,                                       //                               .mem_cas_n
		output wire [0:0]   memory_0_mem_we_n,                                        //                               .mem_we_n
		output wire         memory_0_mem_reset_n,                                     //                               .mem_reset_n
		inout  wire [31:0]  memory_0_mem_dq,                                          //                               .mem_dq
		inout  wire [3:0]   memory_0_mem_dqs,                                         //                               .mem_dqs
		inout  wire [3:0]   memory_0_mem_dqs_n,                                       //                               .mem_dqs_n
		output wire [0:0]   memory_0_mem_odt,                                         //                               .mem_odt
		input  wire         oct_rzqin,                                                //                            oct.rzqin
		output wire         mem_if_ddr3_emif_0_status_local_init_done,                //      mem_if_ddr3_emif_0_status.local_init_done
		output wire         mem_if_ddr3_emif_0_status_local_cal_success,              //                               .local_cal_success
		output wire         mem_if_ddr3_emif_0_status_local_cal_fail,                 //                               .local_cal_fail
		output wire         mem_if_ddr3_emif_0_pll_sharing_pll_mem_clk,               // mem_if_ddr3_emif_0_pll_sharing.pll_mem_clk
		output wire         mem_if_ddr3_emif_0_pll_sharing_pll_write_clk,             //                               .pll_write_clk
		output wire         mem_if_ddr3_emif_0_pll_sharing_pll_locked,                //                               .pll_locked
		output wire         mem_if_ddr3_emif_0_pll_sharing_pll_write_clk_pre_phy_clk, //                               .pll_write_clk_pre_phy_clk
		output wire         mem_if_ddr3_emif_0_pll_sharing_pll_addr_cmd_clk,          //                               .pll_addr_cmd_clk
		output wire         mem_if_ddr3_emif_0_pll_sharing_pll_avl_clk,               //                               .pll_avl_clk
		output wire         mem_if_ddr3_emif_0_pll_sharing_pll_config_clk,            //                               .pll_config_clk
		output wire         mem_if_ddr3_emif_0_pll_sharing_pll_dr_clk,                //                               .pll_dr_clk
		output wire         mem_if_ddr3_emif_0_pll_sharing_pll_dr_clk_pre_phy_clk,    //                               .pll_dr_clk_pre_phy_clk
		output wire         mem_if_ddr3_emif_0_pll_sharing_pll_mem_phy_clk,           //                               .pll_mem_phy_clk
		output wire         mem_if_ddr3_emif_0_pll_sharing_afi_phy_clk,               //                               .afi_phy_clk
		output wire         mem_if_ddr3_emif_0_pll_sharing_pll_avl_phy_clk,           //                               .pll_avl_phy_clk
		output wire         afi_clk_clk,                                              //                        afi_clk.clk
		output wire         mrx_waitrequest,                                          //                            mrx.waitrequest
		output wire [127:0] mrx_readdata,                                             //                               .readdata
		output wire         mrx_readdatavalid,                                        //                               .readdatavalid
		input  wire [5:0]   mrx_burstcount,                                           //                               .burstcount
		input  wire [127:0] mrx_writedata,                                            //                               .writedata
		input  wire [25:0]  mrx_address,                                              //                               .address
		input  wire         mrx_write,                                                //                               .write
		input  wire         mrx_read,                                                 //                               .read
		input  wire [15:0]  mrx_byteenable,                                           //                               .byteenable
		input  wire         mrx_debugaccess,                                          //                               .debugaccess
		output wire         mr0_waitrequest,                                          //                            mr0.waitrequest
		output wire [127:0] mr0_readdata,                                             //                               .readdata
		output wire         mr0_readdatavalid,                                        //                               .readdatavalid
		input  wire [5:0]   mr0_burstcount,                                           //                               .burstcount
		input  wire [127:0] mr0_writedata,                                            //                               .writedata
		input  wire [25:0]  mr0_address,                                              //                               .address
		input  wire         mr0_write,                                                //                               .write
		input  wire         mr0_read,                                                 //                               .read
		input  wire [15:0]  mr0_byteenable,                                           //                               .byteenable
		input  wire         mr0_debugaccess,                                          //                               .debugaccess
		output wire         mr1_waitrequest,                                          //                            mr1.waitrequest
		output wire [127:0] mr1_readdata,                                             //                               .readdata
		output wire         mr1_readdatavalid,                                        //                               .readdatavalid
		input  wire [5:0]   mr1_burstcount,                                           //                               .burstcount
		input  wire [127:0] mr1_writedata,                                            //                               .writedata
		input  wire [25:0]  mr1_address,                                              //                               .address
		input  wire         mr1_write,                                                //                               .write
		input  wire         mr1_read,                                                 //                               .read
		input  wire [15:0]  mr1_byteenable,                                           //                               .byteenable
		input  wire         mr1_debugaccess,                                          //                               .debugaccess
		output wire         mr2_waitrequest,                                          //                            mr2.waitrequest
		output wire [127:0] mr2_readdata,                                             //                               .readdata
		output wire         mr2_readdatavalid,                                        //                               .readdatavalid
		input  wire [5:0]   mr2_burstcount,                                           //                               .burstcount
		input  wire [127:0] mr2_writedata,                                            //                               .writedata
		input  wire [25:0]  mr2_address,                                              //                               .address
		input  wire         mr2_write,                                                //                               .write
		input  wire         mr2_read,                                                 //                               .read
		input  wire [15:0]  mr2_byteenable,                                           //                               .byteenable
		input  wire         mr2_debugaccess,                                          //                               .debugaccess
		output wire         mr3_waitrequest,                                          //                            mr3.waitrequest
		output wire [127:0] mr3_readdata,                                             //                               .readdata
		output wire         mr3_readdatavalid,                                        //                               .readdatavalid
		input  wire [5:0]   mr3_burstcount,                                           //                               .burstcount
		input  wire [127:0] mr3_writedata,                                            //                               .writedata
		input  wire [25:0]  mr3_address,                                              //                               .address
		input  wire         mr3_write,                                                //                               .write
		input  wire         mr3_read,                                                 //                               .read
		input  wire [15:0]  mr3_byteenable,                                           //                               .byteenable
		input  wire         mr3_debugaccess,                                          //                               .debugaccess
		output wire         mwx_waitrequest,                                          //                            mwx.waitrequest
		output wire [127:0] mwx_readdata,                                             //                               .readdata
		output wire         mwx_readdatavalid,                                        //                               .readdatavalid
		input  wire [5:0]   mwx_burstcount,                                           //                               .burstcount
		input  wire [127:0] mwx_writedata,                                            //                               .writedata
		input  wire [25:0]  mwx_address,                                              //                               .address
		input  wire         mwx_write,                                                //                               .write
		input  wire         mwx_read,                                                 //                               .read
		input  wire [15:0]  mwx_byteenable,                                           //                               .byteenable
		input  wire         mwx_debugaccess,                                          //                               .debugaccess
		output wire         mw0_waitrequest,                                          //                            mw0.waitrequest
		output wire [127:0] mw0_readdata,                                             //                               .readdata
		output wire         mw0_readdatavalid,                                        //                               .readdatavalid
		input  wire [5:0]   mw0_burstcount,                                           //                               .burstcount
		input  wire [127:0] mw0_writedata,                                            //                               .writedata
		input  wire [25:0]  mw0_address,                                              //                               .address
		input  wire         mw0_write,                                                //                               .write
		input  wire         mw0_read,                                                 //                               .read
		input  wire [15:0]  mw0_byteenable,                                           //                               .byteenable
		input  wire         mw0_debugaccess,                                          //                               .debugaccess
		output wire         mw1_waitrequest,                                          //                            mw1.waitrequest
		output wire [127:0] mw1_readdata,                                             //                               .readdata
		output wire         mw1_readdatavalid,                                        //                               .readdatavalid
		input  wire [5:0]   mw1_burstcount,                                           //                               .burstcount
		input  wire [127:0] mw1_writedata,                                            //                               .writedata
		input  wire [25:0]  mw1_address,                                              //                               .address
		input  wire         mw1_write,                                                //                               .write
		input  wire         mw1_read,                                                 //                               .read
		input  wire [15:0]  mw1_byteenable,                                           //                               .byteenable
		input  wire         mw1_debugaccess,                                          //                               .debugaccess
		output wire         mw2_waitrequest,                                          //                            mw2.waitrequest
		output wire [127:0] mw2_readdata,                                             //                               .readdata
		output wire         mw2_readdatavalid,                                        //                               .readdatavalid
		input  wire [5:0]   mw2_burstcount,                                           //                               .burstcount
		input  wire [127:0] mw2_writedata,                                            //                               .writedata
		input  wire [25:0]  mw2_address,                                              //                               .address
		input  wire         mw2_write,                                                //                               .write
		input  wire         mw2_read,                                                 //                               .read
		input  wire [15:0]  mw2_byteenable,                                           //                               .byteenable
		input  wire         mw2_debugaccess,                                          //                               .debugaccess
		output wire         mw3_waitrequest,                                          //                            mw3.waitrequest
		output wire [127:0] mw3_readdata,                                             //                               .readdata
		output wire         mw3_readdatavalid,                                        //                               .readdatavalid
		input  wire [5:0]   mw3_burstcount,                                           //                               .burstcount
		input  wire [127:0] mw3_writedata,                                            //                               .writedata
		input  wire [25:0]  mw3_address,                                              //                               .address
		input  wire         mw3_write,                                                //                               .write
		input  wire         mw3_read,                                                 //                               .read
		input  wire [15:0]  mw3_byteenable,                                           //                               .byteenable
		input  wire         mw3_debugaccess,                                          //                               .debugaccess
		output wire         hps_waitrequest,                                          //                            hps.waitrequest
		output wire [127:0] hps_readdata,                                             //                               .readdata
		output wire         hps_readdatavalid,                                        //                               .readdatavalid
		input  wire [5:0]   hps_burstcount,                                           //                               .burstcount
		input  wire [127:0] hps_writedata,                                            //                               .writedata
		input  wire [25:0]  hps_address,                                              //                               .address
		input  wire         hps_write,                                                //                               .write
		input  wire         hps_read,                                                 //                               .read
		input  wire [15:0]  hps_byteenable,                                           //                               .byteenable
		input  wire         hps_debugaccess,                                          //                               .debugaccess
		output wire         mwa_waitrequest,                                          //                            mwa.waitrequest
		output wire [127:0] mwa_readdata,                                             //                               .readdata
		output wire         mwa_readdatavalid,                                        //                               .readdatavalid
		input  wire [5:0]   mwa_burstcount,                                           //                               .burstcount
		input  wire [127:0] mwa_writedata,                                            //                               .writedata
		input  wire [25:0]  mwa_address,                                              //                               .address
		input  wire         mwa_write,                                                //                               .write
		input  wire         mwa_read,                                                 //                               .read
		input  wire [15:0]  mwa_byteenable,                                           //                               .byteenable
		input  wire         mwa_debugaccess,                                          //                               .debugaccess
		input  wire         hps_clk_clk                                               //                        hps_clk.clk
	);

	wire    [5:0] mm_bridge_7_m0_burstcount;                                     // mm_bridge_7:m0_burstcount -> mm_interconnect_0:mm_bridge_7_m0_burstcount
	wire          mm_bridge_7_m0_waitrequest;                                    // mm_interconnect_0:mm_bridge_7_m0_waitrequest -> mm_bridge_7:m0_waitrequest
	wire   [25:0] mm_bridge_7_m0_address;                                        // mm_bridge_7:m0_address -> mm_interconnect_0:mm_bridge_7_m0_address
	wire  [127:0] mm_bridge_7_m0_writedata;                                      // mm_bridge_7:m0_writedata -> mm_interconnect_0:mm_bridge_7_m0_writedata
	wire          mm_bridge_7_m0_write;                                          // mm_bridge_7:m0_write -> mm_interconnect_0:mm_bridge_7_m0_write
	wire          mm_bridge_7_m0_read;                                           // mm_bridge_7:m0_read -> mm_interconnect_0:mm_bridge_7_m0_read
	wire  [127:0] mm_bridge_7_m0_readdata;                                       // mm_interconnect_0:mm_bridge_7_m0_readdata -> mm_bridge_7:m0_readdata
	wire          mm_bridge_7_m0_debugaccess;                                    // mm_bridge_7:m0_debugaccess -> mm_interconnect_0:mm_bridge_7_m0_debugaccess
	wire   [15:0] mm_bridge_7_m0_byteenable;                                     // mm_bridge_7:m0_byteenable -> mm_interconnect_0:mm_bridge_7_m0_byteenable
	wire          mm_bridge_7_m0_readdatavalid;                                  // mm_interconnect_0:mm_bridge_7_m0_readdatavalid -> mm_bridge_7:m0_readdatavalid
	wire    [5:0] mm_bridge_5_m0_burstcount;                                     // mm_bridge_5:m0_burstcount -> mm_interconnect_0:mm_bridge_5_m0_burstcount
	wire          mm_bridge_5_m0_waitrequest;                                    // mm_interconnect_0:mm_bridge_5_m0_waitrequest -> mm_bridge_5:m0_waitrequest
	wire   [25:0] mm_bridge_5_m0_address;                                        // mm_bridge_5:m0_address -> mm_interconnect_0:mm_bridge_5_m0_address
	wire  [127:0] mm_bridge_5_m0_writedata;                                      // mm_bridge_5:m0_writedata -> mm_interconnect_0:mm_bridge_5_m0_writedata
	wire          mm_bridge_5_m0_write;                                          // mm_bridge_5:m0_write -> mm_interconnect_0:mm_bridge_5_m0_write
	wire          mm_bridge_5_m0_read;                                           // mm_bridge_5:m0_read -> mm_interconnect_0:mm_bridge_5_m0_read
	wire  [127:0] mm_bridge_5_m0_readdata;                                       // mm_interconnect_0:mm_bridge_5_m0_readdata -> mm_bridge_5:m0_readdata
	wire          mm_bridge_5_m0_debugaccess;                                    // mm_bridge_5:m0_debugaccess -> mm_interconnect_0:mm_bridge_5_m0_debugaccess
	wire   [15:0] mm_bridge_5_m0_byteenable;                                     // mm_bridge_5:m0_byteenable -> mm_interconnect_0:mm_bridge_5_m0_byteenable
	wire          mm_bridge_5_m0_readdatavalid;                                  // mm_interconnect_0:mm_bridge_5_m0_readdatavalid -> mm_bridge_5:m0_readdatavalid
	wire    [5:0] mm_bridge_0_m0_burstcount;                                     // mm_bridge_0:m0_burstcount -> mm_interconnect_0:mm_bridge_0_m0_burstcount
	wire          mm_bridge_0_m0_waitrequest;                                    // mm_interconnect_0:mm_bridge_0_m0_waitrequest -> mm_bridge_0:m0_waitrequest
	wire   [25:0] mm_bridge_0_m0_address;                                        // mm_bridge_0:m0_address -> mm_interconnect_0:mm_bridge_0_m0_address
	wire  [127:0] mm_bridge_0_m0_writedata;                                      // mm_bridge_0:m0_writedata -> mm_interconnect_0:mm_bridge_0_m0_writedata
	wire          mm_bridge_0_m0_write;                                          // mm_bridge_0:m0_write -> mm_interconnect_0:mm_bridge_0_m0_write
	wire          mm_bridge_0_m0_read;                                           // mm_bridge_0:m0_read -> mm_interconnect_0:mm_bridge_0_m0_read
	wire  [127:0] mm_bridge_0_m0_readdata;                                       // mm_interconnect_0:mm_bridge_0_m0_readdata -> mm_bridge_0:m0_readdata
	wire          mm_bridge_0_m0_debugaccess;                                    // mm_bridge_0:m0_debugaccess -> mm_interconnect_0:mm_bridge_0_m0_debugaccess
	wire   [15:0] mm_bridge_0_m0_byteenable;                                     // mm_bridge_0:m0_byteenable -> mm_interconnect_0:mm_bridge_0_m0_byteenable
	wire          mm_bridge_0_m0_readdatavalid;                                  // mm_interconnect_0:mm_bridge_0_m0_readdatavalid -> mm_bridge_0:m0_readdatavalid
	wire    [5:0] mm_bridge_6_m0_burstcount;                                     // mm_bridge_6:m0_burstcount -> mm_interconnect_0:mm_bridge_6_m0_burstcount
	wire          mm_bridge_6_m0_waitrequest;                                    // mm_interconnect_0:mm_bridge_6_m0_waitrequest -> mm_bridge_6:m0_waitrequest
	wire   [25:0] mm_bridge_6_m0_address;                                        // mm_bridge_6:m0_address -> mm_interconnect_0:mm_bridge_6_m0_address
	wire  [127:0] mm_bridge_6_m0_writedata;                                      // mm_bridge_6:m0_writedata -> mm_interconnect_0:mm_bridge_6_m0_writedata
	wire          mm_bridge_6_m0_write;                                          // mm_bridge_6:m0_write -> mm_interconnect_0:mm_bridge_6_m0_write
	wire          mm_bridge_6_m0_read;                                           // mm_bridge_6:m0_read -> mm_interconnect_0:mm_bridge_6_m0_read
	wire  [127:0] mm_bridge_6_m0_readdata;                                       // mm_interconnect_0:mm_bridge_6_m0_readdata -> mm_bridge_6:m0_readdata
	wire          mm_bridge_6_m0_debugaccess;                                    // mm_bridge_6:m0_debugaccess -> mm_interconnect_0:mm_bridge_6_m0_debugaccess
	wire   [15:0] mm_bridge_6_m0_byteenable;                                     // mm_bridge_6:m0_byteenable -> mm_interconnect_0:mm_bridge_6_m0_byteenable
	wire          mm_bridge_6_m0_readdatavalid;                                  // mm_interconnect_0:mm_bridge_6_m0_readdatavalid -> mm_bridge_6:m0_readdatavalid
	wire    [5:0] mm_bridge_9_m0_burstcount;                                     // mm_bridge_9:m0_burstcount -> mm_interconnect_0:mm_bridge_9_m0_burstcount
	wire          mm_bridge_9_m0_waitrequest;                                    // mm_interconnect_0:mm_bridge_9_m0_waitrequest -> mm_bridge_9:m0_waitrequest
	wire   [25:0] mm_bridge_9_m0_address;                                        // mm_bridge_9:m0_address -> mm_interconnect_0:mm_bridge_9_m0_address
	wire  [127:0] mm_bridge_9_m0_writedata;                                      // mm_bridge_9:m0_writedata -> mm_interconnect_0:mm_bridge_9_m0_writedata
	wire          mm_bridge_9_m0_write;                                          // mm_bridge_9:m0_write -> mm_interconnect_0:mm_bridge_9_m0_write
	wire          mm_bridge_9_m0_read;                                           // mm_bridge_9:m0_read -> mm_interconnect_0:mm_bridge_9_m0_read
	wire  [127:0] mm_bridge_9_m0_readdata;                                       // mm_interconnect_0:mm_bridge_9_m0_readdata -> mm_bridge_9:m0_readdata
	wire          mm_bridge_9_m0_debugaccess;                                    // mm_bridge_9:m0_debugaccess -> mm_interconnect_0:mm_bridge_9_m0_debugaccess
	wire   [15:0] mm_bridge_9_m0_byteenable;                                     // mm_bridge_9:m0_byteenable -> mm_interconnect_0:mm_bridge_9_m0_byteenable
	wire          mm_bridge_9_m0_readdatavalid;                                  // mm_interconnect_0:mm_bridge_9_m0_readdatavalid -> mm_bridge_9:m0_readdatavalid
	wire    [5:0] mm_bridge_11_m0_burstcount;                                    // mm_bridge_11:m0_burstcount -> mm_interconnect_0:mm_bridge_11_m0_burstcount
	wire          mm_bridge_11_m0_waitrequest;                                   // mm_interconnect_0:mm_bridge_11_m0_waitrequest -> mm_bridge_11:m0_waitrequest
	wire   [25:0] mm_bridge_11_m0_address;                                       // mm_bridge_11:m0_address -> mm_interconnect_0:mm_bridge_11_m0_address
	wire  [127:0] mm_bridge_11_m0_writedata;                                     // mm_bridge_11:m0_writedata -> mm_interconnect_0:mm_bridge_11_m0_writedata
	wire          mm_bridge_11_m0_write;                                         // mm_bridge_11:m0_write -> mm_interconnect_0:mm_bridge_11_m0_write
	wire          mm_bridge_11_m0_read;                                          // mm_bridge_11:m0_read -> mm_interconnect_0:mm_bridge_11_m0_read
	wire  [127:0] mm_bridge_11_m0_readdata;                                      // mm_interconnect_0:mm_bridge_11_m0_readdata -> mm_bridge_11:m0_readdata
	wire          mm_bridge_11_m0_debugaccess;                                   // mm_bridge_11:m0_debugaccess -> mm_interconnect_0:mm_bridge_11_m0_debugaccess
	wire   [15:0] mm_bridge_11_m0_byteenable;                                    // mm_bridge_11:m0_byteenable -> mm_interconnect_0:mm_bridge_11_m0_byteenable
	wire          mm_bridge_11_m0_readdatavalid;                                 // mm_interconnect_0:mm_bridge_11_m0_readdatavalid -> mm_bridge_11:m0_readdatavalid
	wire    [5:0] mm_bridge_3_m0_burstcount;                                     // mm_bridge_3:m0_burstcount -> mm_interconnect_0:mm_bridge_3_m0_burstcount
	wire          mm_bridge_3_m0_waitrequest;                                    // mm_interconnect_0:mm_bridge_3_m0_waitrequest -> mm_bridge_3:m0_waitrequest
	wire   [25:0] mm_bridge_3_m0_address;                                        // mm_bridge_3:m0_address -> mm_interconnect_0:mm_bridge_3_m0_address
	wire  [127:0] mm_bridge_3_m0_writedata;                                      // mm_bridge_3:m0_writedata -> mm_interconnect_0:mm_bridge_3_m0_writedata
	wire          mm_bridge_3_m0_write;                                          // mm_bridge_3:m0_write -> mm_interconnect_0:mm_bridge_3_m0_write
	wire          mm_bridge_3_m0_read;                                           // mm_bridge_3:m0_read -> mm_interconnect_0:mm_bridge_3_m0_read
	wire  [127:0] mm_bridge_3_m0_readdata;                                       // mm_interconnect_0:mm_bridge_3_m0_readdata -> mm_bridge_3:m0_readdata
	wire          mm_bridge_3_m0_debugaccess;                                    // mm_bridge_3:m0_debugaccess -> mm_interconnect_0:mm_bridge_3_m0_debugaccess
	wire   [15:0] mm_bridge_3_m0_byteenable;                                     // mm_bridge_3:m0_byteenable -> mm_interconnect_0:mm_bridge_3_m0_byteenable
	wire          mm_bridge_3_m0_readdatavalid;                                  // mm_interconnect_0:mm_bridge_3_m0_readdatavalid -> mm_bridge_3:m0_readdatavalid
	wire    [5:0] mm_bridge_10_m0_burstcount;                                    // mm_bridge_10:m0_burstcount -> mm_interconnect_0:mm_bridge_10_m0_burstcount
	wire          mm_bridge_10_m0_waitrequest;                                   // mm_interconnect_0:mm_bridge_10_m0_waitrequest -> mm_bridge_10:m0_waitrequest
	wire   [25:0] mm_bridge_10_m0_address;                                       // mm_bridge_10:m0_address -> mm_interconnect_0:mm_bridge_10_m0_address
	wire  [127:0] mm_bridge_10_m0_writedata;                                     // mm_bridge_10:m0_writedata -> mm_interconnect_0:mm_bridge_10_m0_writedata
	wire          mm_bridge_10_m0_write;                                         // mm_bridge_10:m0_write -> mm_interconnect_0:mm_bridge_10_m0_write
	wire          mm_bridge_10_m0_read;                                          // mm_bridge_10:m0_read -> mm_interconnect_0:mm_bridge_10_m0_read
	wire  [127:0] mm_bridge_10_m0_readdata;                                      // mm_interconnect_0:mm_bridge_10_m0_readdata -> mm_bridge_10:m0_readdata
	wire          mm_bridge_10_m0_debugaccess;                                   // mm_bridge_10:m0_debugaccess -> mm_interconnect_0:mm_bridge_10_m0_debugaccess
	wire   [15:0] mm_bridge_10_m0_byteenable;                                    // mm_bridge_10:m0_byteenable -> mm_interconnect_0:mm_bridge_10_m0_byteenable
	wire          mm_bridge_10_m0_readdatavalid;                                 // mm_interconnect_0:mm_bridge_10_m0_readdatavalid -> mm_bridge_10:m0_readdatavalid
	wire    [5:0] mm_bridge_2_m0_burstcount;                                     // mm_bridge_2:m0_burstcount -> mm_interconnect_0:mm_bridge_2_m0_burstcount
	wire          mm_bridge_2_m0_waitrequest;                                    // mm_interconnect_0:mm_bridge_2_m0_waitrequest -> mm_bridge_2:m0_waitrequest
	wire   [25:0] mm_bridge_2_m0_address;                                        // mm_bridge_2:m0_address -> mm_interconnect_0:mm_bridge_2_m0_address
	wire  [127:0] mm_bridge_2_m0_writedata;                                      // mm_bridge_2:m0_writedata -> mm_interconnect_0:mm_bridge_2_m0_writedata
	wire          mm_bridge_2_m0_write;                                          // mm_bridge_2:m0_write -> mm_interconnect_0:mm_bridge_2_m0_write
	wire          mm_bridge_2_m0_read;                                           // mm_bridge_2:m0_read -> mm_interconnect_0:mm_bridge_2_m0_read
	wire  [127:0] mm_bridge_2_m0_readdata;                                       // mm_interconnect_0:mm_bridge_2_m0_readdata -> mm_bridge_2:m0_readdata
	wire          mm_bridge_2_m0_debugaccess;                                    // mm_bridge_2:m0_debugaccess -> mm_interconnect_0:mm_bridge_2_m0_debugaccess
	wire   [15:0] mm_bridge_2_m0_byteenable;                                     // mm_bridge_2:m0_byteenable -> mm_interconnect_0:mm_bridge_2_m0_byteenable
	wire          mm_bridge_2_m0_readdatavalid;                                  // mm_interconnect_0:mm_bridge_2_m0_readdatavalid -> mm_bridge_2:m0_readdatavalid
	wire    [5:0] mm_bridge_1_m0_burstcount;                                     // mm_bridge_1:m0_burstcount -> mm_interconnect_0:mm_bridge_1_m0_burstcount
	wire          mm_bridge_1_m0_waitrequest;                                    // mm_interconnect_0:mm_bridge_1_m0_waitrequest -> mm_bridge_1:m0_waitrequest
	wire   [25:0] mm_bridge_1_m0_address;                                        // mm_bridge_1:m0_address -> mm_interconnect_0:mm_bridge_1_m0_address
	wire  [127:0] mm_bridge_1_m0_writedata;                                      // mm_bridge_1:m0_writedata -> mm_interconnect_0:mm_bridge_1_m0_writedata
	wire          mm_bridge_1_m0_write;                                          // mm_bridge_1:m0_write -> mm_interconnect_0:mm_bridge_1_m0_write
	wire          mm_bridge_1_m0_read;                                           // mm_bridge_1:m0_read -> mm_interconnect_0:mm_bridge_1_m0_read
	wire  [127:0] mm_bridge_1_m0_readdata;                                       // mm_interconnect_0:mm_bridge_1_m0_readdata -> mm_bridge_1:m0_readdata
	wire          mm_bridge_1_m0_debugaccess;                                    // mm_bridge_1:m0_debugaccess -> mm_interconnect_0:mm_bridge_1_m0_debugaccess
	wire   [15:0] mm_bridge_1_m0_byteenable;                                     // mm_bridge_1:m0_byteenable -> mm_interconnect_0:mm_bridge_1_m0_byteenable
	wire          mm_bridge_1_m0_readdatavalid;                                  // mm_interconnect_0:mm_bridge_1_m0_readdatavalid -> mm_bridge_1:m0_readdatavalid
	wire    [5:0] mm_bridge_8_m0_burstcount;                                     // mm_bridge_8:m0_burstcount -> mm_interconnect_0:mm_bridge_8_m0_burstcount
	wire          mm_bridge_8_m0_waitrequest;                                    // mm_interconnect_0:mm_bridge_8_m0_waitrequest -> mm_bridge_8:m0_waitrequest
	wire   [25:0] mm_bridge_8_m0_address;                                        // mm_bridge_8:m0_address -> mm_interconnect_0:mm_bridge_8_m0_address
	wire  [127:0] mm_bridge_8_m0_writedata;                                      // mm_bridge_8:m0_writedata -> mm_interconnect_0:mm_bridge_8_m0_writedata
	wire          mm_bridge_8_m0_write;                                          // mm_bridge_8:m0_write -> mm_interconnect_0:mm_bridge_8_m0_write
	wire          mm_bridge_8_m0_read;                                           // mm_bridge_8:m0_read -> mm_interconnect_0:mm_bridge_8_m0_read
	wire  [127:0] mm_bridge_8_m0_readdata;                                       // mm_interconnect_0:mm_bridge_8_m0_readdata -> mm_bridge_8:m0_readdata
	wire          mm_bridge_8_m0_debugaccess;                                    // mm_bridge_8:m0_debugaccess -> mm_interconnect_0:mm_bridge_8_m0_debugaccess
	wire   [15:0] mm_bridge_8_m0_byteenable;                                     // mm_bridge_8:m0_byteenable -> mm_interconnect_0:mm_bridge_8_m0_byteenable
	wire          mm_bridge_8_m0_readdatavalid;                                  // mm_interconnect_0:mm_bridge_8_m0_readdatavalid -> mm_bridge_8:m0_readdatavalid
	wire          mm_interconnect_0_mem_if_ddr3_emif_0_avl_0_waitrequest;        // mem_if_ddr3_emif_0:avl_ready_0 -> mm_interconnect_0:mem_if_ddr3_emif_0_avl_0_waitrequest
	wire    [5:0] mm_interconnect_0_mem_if_ddr3_emif_0_avl_0_burstcount;         // mm_interconnect_0:mem_if_ddr3_emif_0_avl_0_burstcount -> mem_if_ddr3_emif_0:avl_size_0
	wire  [127:0] mm_interconnect_0_mem_if_ddr3_emif_0_avl_0_writedata;          // mm_interconnect_0:mem_if_ddr3_emif_0_avl_0_writedata -> mem_if_ddr3_emif_0:avl_wdata_0
	wire   [25:0] mm_interconnect_0_mem_if_ddr3_emif_0_avl_0_address;            // mm_interconnect_0:mem_if_ddr3_emif_0_avl_0_address -> mem_if_ddr3_emif_0:avl_addr_0
	wire          mm_interconnect_0_mem_if_ddr3_emif_0_avl_0_write;              // mm_interconnect_0:mem_if_ddr3_emif_0_avl_0_write -> mem_if_ddr3_emif_0:avl_write_req_0
	wire          mm_interconnect_0_mem_if_ddr3_emif_0_avl_0_beginbursttransfer; // mm_interconnect_0:mem_if_ddr3_emif_0_avl_0_beginbursttransfer -> mem_if_ddr3_emif_0:avl_burstbegin_0
	wire          mm_interconnect_0_mem_if_ddr3_emif_0_avl_0_read;               // mm_interconnect_0:mem_if_ddr3_emif_0_avl_0_read -> mem_if_ddr3_emif_0:avl_read_req_0
	wire  [127:0] mm_interconnect_0_mem_if_ddr3_emif_0_avl_0_readdata;           // mem_if_ddr3_emif_0:avl_rdata_0 -> mm_interconnect_0:mem_if_ddr3_emif_0_avl_0_readdata
	wire          mm_interconnect_0_mem_if_ddr3_emif_0_avl_0_readdatavalid;      // mem_if_ddr3_emif_0:avl_rdata_valid_0 -> mm_interconnect_0:mem_if_ddr3_emif_0_avl_0_readdatavalid
	wire   [15:0] mm_interconnect_0_mem_if_ddr3_emif_0_avl_0_byteenable;         // mm_interconnect_0:mem_if_ddr3_emif_0_avl_0_byteenable -> mem_if_ddr3_emif_0:avl_be_0
	wire    [5:0] mm_bridge_4_m0_burstcount;                                     // mm_bridge_4:m0_burstcount -> mm_interconnect_0:mm_bridge_4_m0_burstcount
	wire          mm_bridge_4_m0_waitrequest;                                    // mm_interconnect_0:mm_bridge_4_m0_waitrequest -> mm_bridge_4:m0_waitrequest
	wire   [25:0] mm_bridge_4_m0_address;                                        // mm_bridge_4:m0_address -> mm_interconnect_0:mm_bridge_4_m0_address
	wire  [127:0] mm_bridge_4_m0_writedata;                                      // mm_bridge_4:m0_writedata -> mm_interconnect_0:mm_bridge_4_m0_writedata
	wire          mm_bridge_4_m0_write;                                          // mm_bridge_4:m0_write -> mm_interconnect_0:mm_bridge_4_m0_write
	wire          mm_bridge_4_m0_read;                                           // mm_bridge_4:m0_read -> mm_interconnect_0:mm_bridge_4_m0_read
	wire  [127:0] mm_bridge_4_m0_readdata;                                       // mm_interconnect_0:mm_bridge_4_m0_readdata -> mm_bridge_4:m0_readdata
	wire          mm_bridge_4_m0_debugaccess;                                    // mm_bridge_4:m0_debugaccess -> mm_interconnect_0:mm_bridge_4_m0_debugaccess
	wire   [15:0] mm_bridge_4_m0_byteenable;                                     // mm_bridge_4:m0_byteenable -> mm_interconnect_0:mm_bridge_4_m0_byteenable
	wire          mm_bridge_4_m0_readdatavalid;                                  // mm_interconnect_0:mm_bridge_4_m0_readdatavalid -> mm_bridge_4:m0_readdatavalid
	wire          rst_controller_reset_out_reset;                                // rst_controller:reset_out -> [mm_bridge_0:reset, mm_bridge_11:reset, mm_bridge_1:reset, mm_bridge_2:reset, mm_bridge_3:reset, mm_bridge_4:reset, mm_bridge_5:reset, mm_bridge_6:reset, mm_bridge_7:reset, mm_bridge_8:reset, mm_bridge_9:reset, mm_interconnect_0:mem_if_ddr3_emif_0_mp_cmd_reset_n_0_reset_bridge_in_reset_reset, mm_interconnect_0:mm_bridge_11_reset_reset_bridge_in_reset_reset]
	wire          rst_controller_001_reset_out_reset;                            // rst_controller_001:reset_out -> [mm_bridge_10:reset, mm_interconnect_0:mm_bridge_10_reset_reset_bridge_in_reset_reset]

	fpga_mem_mem_if_ddr3_emif_0 mem_if_ddr3_emif_0 (
		.pll_ref_clk                (clk_clk),                                                       //        pll_ref_clk.clk
		.global_reset_n             (reset_reset_n),                                                 //       global_reset.reset_n
		.soft_reset_n               (reset_reset_n),                                                 //         soft_reset.reset_n
		.afi_clk                    (),                                                              //            afi_clk.clk
		.afi_half_clk               (afi_clk_clk),                                                   //       afi_half_clk.clk
		.afi_reset_n                (),                                                              //          afi_reset.reset_n
		.afi_reset_export_n         (),                                                              //   afi_reset_export.reset_n
		.mem_a                      (memory_0_mem_a),                                                //             memory.mem_a
		.mem_ba                     (memory_0_mem_ba),                                               //                   .mem_ba
		.mem_ck                     (memory_0_mem_ck),                                               //                   .mem_ck
		.mem_ck_n                   (memory_0_mem_ck_n),                                             //                   .mem_ck_n
		.mem_cke                    (memory_0_mem_cke),                                              //                   .mem_cke
		.mem_cs_n                   (memory_0_mem_cs_n),                                             //                   .mem_cs_n
		.mem_dm                     (memory_0_mem_dm),                                               //                   .mem_dm
		.mem_ras_n                  (memory_0_mem_ras_n),                                            //                   .mem_ras_n
		.mem_cas_n                  (memory_0_mem_cas_n),                                            //                   .mem_cas_n
		.mem_we_n                   (memory_0_mem_we_n),                                             //                   .mem_we_n
		.mem_reset_n                (memory_0_mem_reset_n),                                          //                   .mem_reset_n
		.mem_dq                     (memory_0_mem_dq),                                               //                   .mem_dq
		.mem_dqs                    (memory_0_mem_dqs),                                              //                   .mem_dqs
		.mem_dqs_n                  (memory_0_mem_dqs_n),                                            //                   .mem_dqs_n
		.mem_odt                    (memory_0_mem_odt),                                              //                   .mem_odt
		.avl_ready_0                (mm_interconnect_0_mem_if_ddr3_emif_0_avl_0_waitrequest),        //              avl_0.waitrequest_n
		.avl_burstbegin_0           (mm_interconnect_0_mem_if_ddr3_emif_0_avl_0_beginbursttransfer), //                   .beginbursttransfer
		.avl_addr_0                 (mm_interconnect_0_mem_if_ddr3_emif_0_avl_0_address),            //                   .address
		.avl_rdata_valid_0          (mm_interconnect_0_mem_if_ddr3_emif_0_avl_0_readdatavalid),      //                   .readdatavalid
		.avl_rdata_0                (mm_interconnect_0_mem_if_ddr3_emif_0_avl_0_readdata),           //                   .readdata
		.avl_wdata_0                (mm_interconnect_0_mem_if_ddr3_emif_0_avl_0_writedata),          //                   .writedata
		.avl_be_0                   (mm_interconnect_0_mem_if_ddr3_emif_0_avl_0_byteenable),         //                   .byteenable
		.avl_read_req_0             (mm_interconnect_0_mem_if_ddr3_emif_0_avl_0_read),               //                   .read
		.avl_write_req_0            (mm_interconnect_0_mem_if_ddr3_emif_0_avl_0_write),              //                   .write
		.avl_size_0                 (mm_interconnect_0_mem_if_ddr3_emif_0_avl_0_burstcount),         //                   .burstcount
		.mp_cmd_clk_0_clk           (afi_clk_clk),                                                   //       mp_cmd_clk_0.clk
		.mp_cmd_reset_n_0_reset_n   (reset_reset_n),                                                 //   mp_cmd_reset_n_0.reset_n
		.mp_rfifo_clk_0_clk         (afi_clk_clk),                                                   //     mp_rfifo_clk_0.clk
		.mp_rfifo_reset_n_0_reset_n (reset_reset_n),                                                 // mp_rfifo_reset_n_0.reset_n
		.mp_wfifo_clk_0_clk         (afi_clk_clk),                                                   //     mp_wfifo_clk_0.clk
		.mp_wfifo_reset_n_0_reset_n (reset_reset_n),                                                 // mp_wfifo_reset_n_0.reset_n
		.mp_rfifo_clk_1_clk         (afi_clk_clk),                                                   //     mp_rfifo_clk_1.clk
		.mp_rfifo_reset_n_1_reset_n (reset_reset_n),                                                 // mp_rfifo_reset_n_1.reset_n
		.mp_wfifo_clk_1_clk         (afi_clk_clk),                                                   //     mp_wfifo_clk_1.clk
		.mp_wfifo_reset_n_1_reset_n (reset_reset_n),                                                 // mp_wfifo_reset_n_1.reset_n
		.local_init_done            (mem_if_ddr3_emif_0_status_local_init_done),                     //             status.local_init_done
		.local_cal_success          (mem_if_ddr3_emif_0_status_local_cal_success),                   //                   .local_cal_success
		.local_cal_fail             (mem_if_ddr3_emif_0_status_local_cal_fail),                      //                   .local_cal_fail
		.oct_rzqin                  (oct_rzqin),                                                     //                oct.rzqin
		.pll_mem_clk                (mem_if_ddr3_emif_0_pll_sharing_pll_mem_clk),                    //        pll_sharing.pll_mem_clk
		.pll_write_clk              (mem_if_ddr3_emif_0_pll_sharing_pll_write_clk),                  //                   .pll_write_clk
		.pll_locked                 (mem_if_ddr3_emif_0_pll_sharing_pll_locked),                     //                   .pll_locked
		.pll_write_clk_pre_phy_clk  (mem_if_ddr3_emif_0_pll_sharing_pll_write_clk_pre_phy_clk),      //                   .pll_write_clk_pre_phy_clk
		.pll_addr_cmd_clk           (mem_if_ddr3_emif_0_pll_sharing_pll_addr_cmd_clk),               //                   .pll_addr_cmd_clk
		.pll_avl_clk                (mem_if_ddr3_emif_0_pll_sharing_pll_avl_clk),                    //                   .pll_avl_clk
		.pll_config_clk             (mem_if_ddr3_emif_0_pll_sharing_pll_config_clk),                 //                   .pll_config_clk
		.pll_dr_clk                 (mem_if_ddr3_emif_0_pll_sharing_pll_dr_clk),                     //                   .pll_dr_clk
		.pll_dr_clk_pre_phy_clk     (mem_if_ddr3_emif_0_pll_sharing_pll_dr_clk_pre_phy_clk),         //                   .pll_dr_clk_pre_phy_clk
		.pll_mem_phy_clk            (mem_if_ddr3_emif_0_pll_sharing_pll_mem_phy_clk),                //                   .pll_mem_phy_clk
		.afi_phy_clk                (mem_if_ddr3_emif_0_pll_sharing_afi_phy_clk),                    //                   .afi_phy_clk
		.pll_avl_phy_clk            (mem_if_ddr3_emif_0_pll_sharing_pll_avl_phy_clk)                 //                   .pll_avl_phy_clk
	);

	altera_avalon_mm_bridge #(
		.DATA_WIDTH        (128),
		.SYMBOL_WIDTH      (8),
		.ADDRESS_WIDTH     (26),
		.BURSTCOUNT_WIDTH  (6),
		.PIPELINE_COMMAND  (1),
		.PIPELINE_RESPONSE (1)
	) mm_bridge_0 (
		.clk              (afi_clk_clk),                    //   clk.clk
		.reset            (rst_controller_reset_out_reset), // reset.reset
		.s0_waitrequest   (mrx_waitrequest),                //    s0.waitrequest
		.s0_readdata      (mrx_readdata),                   //      .readdata
		.s0_readdatavalid (mrx_readdatavalid),              //      .readdatavalid
		.s0_burstcount    (mrx_burstcount),                 //      .burstcount
		.s0_writedata     (mrx_writedata),                  //      .writedata
		.s0_address       (mrx_address),                    //      .address
		.s0_write         (mrx_write),                      //      .write
		.s0_read          (mrx_read),                       //      .read
		.s0_byteenable    (mrx_byteenable),                 //      .byteenable
		.s0_debugaccess   (mrx_debugaccess),                //      .debugaccess
		.m0_waitrequest   (mm_bridge_0_m0_waitrequest),     //    m0.waitrequest
		.m0_readdata      (mm_bridge_0_m0_readdata),        //      .readdata
		.m0_readdatavalid (mm_bridge_0_m0_readdatavalid),   //      .readdatavalid
		.m0_burstcount    (mm_bridge_0_m0_burstcount),      //      .burstcount
		.m0_writedata     (mm_bridge_0_m0_writedata),       //      .writedata
		.m0_address       (mm_bridge_0_m0_address),         //      .address
		.m0_write         (mm_bridge_0_m0_write),           //      .write
		.m0_read          (mm_bridge_0_m0_read),            //      .read
		.m0_byteenable    (mm_bridge_0_m0_byteenable),      //      .byteenable
		.m0_debugaccess   (mm_bridge_0_m0_debugaccess)      //      .debugaccess
	);

	altera_avalon_mm_bridge #(
		.DATA_WIDTH        (128),
		.SYMBOL_WIDTH      (8),
		.ADDRESS_WIDTH     (26),
		.BURSTCOUNT_WIDTH  (6),
		.PIPELINE_COMMAND  (1),
		.PIPELINE_RESPONSE (1)
	) mm_bridge_1 (
		.clk              (afi_clk_clk),                    //   clk.clk
		.reset            (rst_controller_reset_out_reset), // reset.reset
		.s0_waitrequest   (mr0_waitrequest),                //    s0.waitrequest
		.s0_readdata      (mr0_readdata),                   //      .readdata
		.s0_readdatavalid (mr0_readdatavalid),              //      .readdatavalid
		.s0_burstcount    (mr0_burstcount),                 //      .burstcount
		.s0_writedata     (mr0_writedata),                  //      .writedata
		.s0_address       (mr0_address),                    //      .address
		.s0_write         (mr0_write),                      //      .write
		.s0_read          (mr0_read),                       //      .read
		.s0_byteenable    (mr0_byteenable),                 //      .byteenable
		.s0_debugaccess   (mr0_debugaccess),                //      .debugaccess
		.m0_waitrequest   (mm_bridge_1_m0_waitrequest),     //    m0.waitrequest
		.m0_readdata      (mm_bridge_1_m0_readdata),        //      .readdata
		.m0_readdatavalid (mm_bridge_1_m0_readdatavalid),   //      .readdatavalid
		.m0_burstcount    (mm_bridge_1_m0_burstcount),      //      .burstcount
		.m0_writedata     (mm_bridge_1_m0_writedata),       //      .writedata
		.m0_address       (mm_bridge_1_m0_address),         //      .address
		.m0_write         (mm_bridge_1_m0_write),           //      .write
		.m0_read          (mm_bridge_1_m0_read),            //      .read
		.m0_byteenable    (mm_bridge_1_m0_byteenable),      //      .byteenable
		.m0_debugaccess   (mm_bridge_1_m0_debugaccess)      //      .debugaccess
	);

	altera_avalon_mm_bridge #(
		.DATA_WIDTH        (128),
		.SYMBOL_WIDTH      (8),
		.ADDRESS_WIDTH     (26),
		.BURSTCOUNT_WIDTH  (6),
		.PIPELINE_COMMAND  (1),
		.PIPELINE_RESPONSE (1)
	) mm_bridge_2 (
		.clk              (afi_clk_clk),                    //   clk.clk
		.reset            (rst_controller_reset_out_reset), // reset.reset
		.s0_waitrequest   (mr1_waitrequest),                //    s0.waitrequest
		.s0_readdata      (mr1_readdata),                   //      .readdata
		.s0_readdatavalid (mr1_readdatavalid),              //      .readdatavalid
		.s0_burstcount    (mr1_burstcount),                 //      .burstcount
		.s0_writedata     (mr1_writedata),                  //      .writedata
		.s0_address       (mr1_address),                    //      .address
		.s0_write         (mr1_write),                      //      .write
		.s0_read          (mr1_read),                       //      .read
		.s0_byteenable    (mr1_byteenable),                 //      .byteenable
		.s0_debugaccess   (mr1_debugaccess),                //      .debugaccess
		.m0_waitrequest   (mm_bridge_2_m0_waitrequest),     //    m0.waitrequest
		.m0_readdata      (mm_bridge_2_m0_readdata),        //      .readdata
		.m0_readdatavalid (mm_bridge_2_m0_readdatavalid),   //      .readdatavalid
		.m0_burstcount    (mm_bridge_2_m0_burstcount),      //      .burstcount
		.m0_writedata     (mm_bridge_2_m0_writedata),       //      .writedata
		.m0_address       (mm_bridge_2_m0_address),         //      .address
		.m0_write         (mm_bridge_2_m0_write),           //      .write
		.m0_read          (mm_bridge_2_m0_read),            //      .read
		.m0_byteenable    (mm_bridge_2_m0_byteenable),      //      .byteenable
		.m0_debugaccess   (mm_bridge_2_m0_debugaccess)      //      .debugaccess
	);

	altera_avalon_mm_bridge #(
		.DATA_WIDTH        (128),
		.SYMBOL_WIDTH      (8),
		.ADDRESS_WIDTH     (26),
		.BURSTCOUNT_WIDTH  (6),
		.PIPELINE_COMMAND  (1),
		.PIPELINE_RESPONSE (1)
	) mm_bridge_3 (
		.clk              (afi_clk_clk),                    //   clk.clk
		.reset            (rst_controller_reset_out_reset), // reset.reset
		.s0_waitrequest   (mr2_waitrequest),                //    s0.waitrequest
		.s0_readdata      (mr2_readdata),                   //      .readdata
		.s0_readdatavalid (mr2_readdatavalid),              //      .readdatavalid
		.s0_burstcount    (mr2_burstcount),                 //      .burstcount
		.s0_writedata     (mr2_writedata),                  //      .writedata
		.s0_address       (mr2_address),                    //      .address
		.s0_write         (mr2_write),                      //      .write
		.s0_read          (mr2_read),                       //      .read
		.s0_byteenable    (mr2_byteenable),                 //      .byteenable
		.s0_debugaccess   (mr2_debugaccess),                //      .debugaccess
		.m0_waitrequest   (mm_bridge_3_m0_waitrequest),     //    m0.waitrequest
		.m0_readdata      (mm_bridge_3_m0_readdata),        //      .readdata
		.m0_readdatavalid (mm_bridge_3_m0_readdatavalid),   //      .readdatavalid
		.m0_burstcount    (mm_bridge_3_m0_burstcount),      //      .burstcount
		.m0_writedata     (mm_bridge_3_m0_writedata),       //      .writedata
		.m0_address       (mm_bridge_3_m0_address),         //      .address
		.m0_write         (mm_bridge_3_m0_write),           //      .write
		.m0_read          (mm_bridge_3_m0_read),            //      .read
		.m0_byteenable    (mm_bridge_3_m0_byteenable),      //      .byteenable
		.m0_debugaccess   (mm_bridge_3_m0_debugaccess)      //      .debugaccess
	);

	altera_avalon_mm_bridge #(
		.DATA_WIDTH        (128),
		.SYMBOL_WIDTH      (8),
		.ADDRESS_WIDTH     (26),
		.BURSTCOUNT_WIDTH  (6),
		.PIPELINE_COMMAND  (1),
		.PIPELINE_RESPONSE (1)
	) mm_bridge_4 (
		.clk              (afi_clk_clk),                    //   clk.clk
		.reset            (rst_controller_reset_out_reset), // reset.reset
		.s0_waitrequest   (mr3_waitrequest),                //    s0.waitrequest
		.s0_readdata      (mr3_readdata),                   //      .readdata
		.s0_readdatavalid (mr3_readdatavalid),              //      .readdatavalid
		.s0_burstcount    (mr3_burstcount),                 //      .burstcount
		.s0_writedata     (mr3_writedata),                  //      .writedata
		.s0_address       (mr3_address),                    //      .address
		.s0_write         (mr3_write),                      //      .write
		.s0_read          (mr3_read),                       //      .read
		.s0_byteenable    (mr3_byteenable),                 //      .byteenable
		.s0_debugaccess   (mr3_debugaccess),                //      .debugaccess
		.m0_waitrequest   (mm_bridge_4_m0_waitrequest),     //    m0.waitrequest
		.m0_readdata      (mm_bridge_4_m0_readdata),        //      .readdata
		.m0_readdatavalid (mm_bridge_4_m0_readdatavalid),   //      .readdatavalid
		.m0_burstcount    (mm_bridge_4_m0_burstcount),      //      .burstcount
		.m0_writedata     (mm_bridge_4_m0_writedata),       //      .writedata
		.m0_address       (mm_bridge_4_m0_address),         //      .address
		.m0_write         (mm_bridge_4_m0_write),           //      .write
		.m0_read          (mm_bridge_4_m0_read),            //      .read
		.m0_byteenable    (mm_bridge_4_m0_byteenable),      //      .byteenable
		.m0_debugaccess   (mm_bridge_4_m0_debugaccess)      //      .debugaccess
	);

	altera_avalon_mm_bridge #(
		.DATA_WIDTH        (128),
		.SYMBOL_WIDTH      (8),
		.ADDRESS_WIDTH     (26),
		.BURSTCOUNT_WIDTH  (6),
		.PIPELINE_COMMAND  (1),
		.PIPELINE_RESPONSE (1)
	) mm_bridge_5 (
		.clk              (afi_clk_clk),                    //   clk.clk
		.reset            (rst_controller_reset_out_reset), // reset.reset
		.s0_waitrequest   (mwx_waitrequest),                //    s0.waitrequest
		.s0_readdata      (mwx_readdata),                   //      .readdata
		.s0_readdatavalid (mwx_readdatavalid),              //      .readdatavalid
		.s0_burstcount    (mwx_burstcount),                 //      .burstcount
		.s0_writedata     (mwx_writedata),                  //      .writedata
		.s0_address       (mwx_address),                    //      .address
		.s0_write         (mwx_write),                      //      .write
		.s0_read          (mwx_read),                       //      .read
		.s0_byteenable    (mwx_byteenable),                 //      .byteenable
		.s0_debugaccess   (mwx_debugaccess),                //      .debugaccess
		.m0_waitrequest   (mm_bridge_5_m0_waitrequest),     //    m0.waitrequest
		.m0_readdata      (mm_bridge_5_m0_readdata),        //      .readdata
		.m0_readdatavalid (mm_bridge_5_m0_readdatavalid),   //      .readdatavalid
		.m0_burstcount    (mm_bridge_5_m0_burstcount),      //      .burstcount
		.m0_writedata     (mm_bridge_5_m0_writedata),       //      .writedata
		.m0_address       (mm_bridge_5_m0_address),         //      .address
		.m0_write         (mm_bridge_5_m0_write),           //      .write
		.m0_read          (mm_bridge_5_m0_read),            //      .read
		.m0_byteenable    (mm_bridge_5_m0_byteenable),      //      .byteenable
		.m0_debugaccess   (mm_bridge_5_m0_debugaccess)      //      .debugaccess
	);

	altera_avalon_mm_bridge #(
		.DATA_WIDTH        (128),
		.SYMBOL_WIDTH      (8),
		.ADDRESS_WIDTH     (26),
		.BURSTCOUNT_WIDTH  (6),
		.PIPELINE_COMMAND  (1),
		.PIPELINE_RESPONSE (1)
	) mm_bridge_6 (
		.clk              (afi_clk_clk),                    //   clk.clk
		.reset            (rst_controller_reset_out_reset), // reset.reset
		.s0_waitrequest   (mw0_waitrequest),                //    s0.waitrequest
		.s0_readdata      (mw0_readdata),                   //      .readdata
		.s0_readdatavalid (mw0_readdatavalid),              //      .readdatavalid
		.s0_burstcount    (mw0_burstcount),                 //      .burstcount
		.s0_writedata     (mw0_writedata),                  //      .writedata
		.s0_address       (mw0_address),                    //      .address
		.s0_write         (mw0_write),                      //      .write
		.s0_read          (mw0_read),                       //      .read
		.s0_byteenable    (mw0_byteenable),                 //      .byteenable
		.s0_debugaccess   (mw0_debugaccess),                //      .debugaccess
		.m0_waitrequest   (mm_bridge_6_m0_waitrequest),     //    m0.waitrequest
		.m0_readdata      (mm_bridge_6_m0_readdata),        //      .readdata
		.m0_readdatavalid (mm_bridge_6_m0_readdatavalid),   //      .readdatavalid
		.m0_burstcount    (mm_bridge_6_m0_burstcount),      //      .burstcount
		.m0_writedata     (mm_bridge_6_m0_writedata),       //      .writedata
		.m0_address       (mm_bridge_6_m0_address),         //      .address
		.m0_write         (mm_bridge_6_m0_write),           //      .write
		.m0_read          (mm_bridge_6_m0_read),            //      .read
		.m0_byteenable    (mm_bridge_6_m0_byteenable),      //      .byteenable
		.m0_debugaccess   (mm_bridge_6_m0_debugaccess)      //      .debugaccess
	);

	altera_avalon_mm_bridge #(
		.DATA_WIDTH        (128),
		.SYMBOL_WIDTH      (8),
		.ADDRESS_WIDTH     (26),
		.BURSTCOUNT_WIDTH  (6),
		.PIPELINE_COMMAND  (1),
		.PIPELINE_RESPONSE (1)
	) mm_bridge_7 (
		.clk              (afi_clk_clk),                    //   clk.clk
		.reset            (rst_controller_reset_out_reset), // reset.reset
		.s0_waitrequest   (mw1_waitrequest),                //    s0.waitrequest
		.s0_readdata      (mw1_readdata),                   //      .readdata
		.s0_readdatavalid (mw1_readdatavalid),              //      .readdatavalid
		.s0_burstcount    (mw1_burstcount),                 //      .burstcount
		.s0_writedata     (mw1_writedata),                  //      .writedata
		.s0_address       (mw1_address),                    //      .address
		.s0_write         (mw1_write),                      //      .write
		.s0_read          (mw1_read),                       //      .read
		.s0_byteenable    (mw1_byteenable),                 //      .byteenable
		.s0_debugaccess   (mw1_debugaccess),                //      .debugaccess
		.m0_waitrequest   (mm_bridge_7_m0_waitrequest),     //    m0.waitrequest
		.m0_readdata      (mm_bridge_7_m0_readdata),        //      .readdata
		.m0_readdatavalid (mm_bridge_7_m0_readdatavalid),   //      .readdatavalid
		.m0_burstcount    (mm_bridge_7_m0_burstcount),      //      .burstcount
		.m0_writedata     (mm_bridge_7_m0_writedata),       //      .writedata
		.m0_address       (mm_bridge_7_m0_address),         //      .address
		.m0_write         (mm_bridge_7_m0_write),           //      .write
		.m0_read          (mm_bridge_7_m0_read),            //      .read
		.m0_byteenable    (mm_bridge_7_m0_byteenable),      //      .byteenable
		.m0_debugaccess   (mm_bridge_7_m0_debugaccess)      //      .debugaccess
	);

	altera_avalon_mm_bridge #(
		.DATA_WIDTH        (128),
		.SYMBOL_WIDTH      (8),
		.ADDRESS_WIDTH     (26),
		.BURSTCOUNT_WIDTH  (6),
		.PIPELINE_COMMAND  (1),
		.PIPELINE_RESPONSE (1)
	) mm_bridge_8 (
		.clk              (afi_clk_clk),                    //   clk.clk
		.reset            (rst_controller_reset_out_reset), // reset.reset
		.s0_waitrequest   (mw2_waitrequest),                //    s0.waitrequest
		.s0_readdata      (mw2_readdata),                   //      .readdata
		.s0_readdatavalid (mw2_readdatavalid),              //      .readdatavalid
		.s0_burstcount    (mw2_burstcount),                 //      .burstcount
		.s0_writedata     (mw2_writedata),                  //      .writedata
		.s0_address       (mw2_address),                    //      .address
		.s0_write         (mw2_write),                      //      .write
		.s0_read          (mw2_read),                       //      .read
		.s0_byteenable    (mw2_byteenable),                 //      .byteenable
		.s0_debugaccess   (mw2_debugaccess),                //      .debugaccess
		.m0_waitrequest   (mm_bridge_8_m0_waitrequest),     //    m0.waitrequest
		.m0_readdata      (mm_bridge_8_m0_readdata),        //      .readdata
		.m0_readdatavalid (mm_bridge_8_m0_readdatavalid),   //      .readdatavalid
		.m0_burstcount    (mm_bridge_8_m0_burstcount),      //      .burstcount
		.m0_writedata     (mm_bridge_8_m0_writedata),       //      .writedata
		.m0_address       (mm_bridge_8_m0_address),         //      .address
		.m0_write         (mm_bridge_8_m0_write),           //      .write
		.m0_read          (mm_bridge_8_m0_read),            //      .read
		.m0_byteenable    (mm_bridge_8_m0_byteenable),      //      .byteenable
		.m0_debugaccess   (mm_bridge_8_m0_debugaccess)      //      .debugaccess
	);

	altera_avalon_mm_bridge #(
		.DATA_WIDTH        (128),
		.SYMBOL_WIDTH      (8),
		.ADDRESS_WIDTH     (26),
		.BURSTCOUNT_WIDTH  (6),
		.PIPELINE_COMMAND  (1),
		.PIPELINE_RESPONSE (1)
	) mm_bridge_9 (
		.clk              (afi_clk_clk),                    //   clk.clk
		.reset            (rst_controller_reset_out_reset), // reset.reset
		.s0_waitrequest   (mw3_waitrequest),                //    s0.waitrequest
		.s0_readdata      (mw3_readdata),                   //      .readdata
		.s0_readdatavalid (mw3_readdatavalid),              //      .readdatavalid
		.s0_burstcount    (mw3_burstcount),                 //      .burstcount
		.s0_writedata     (mw3_writedata),                  //      .writedata
		.s0_address       (mw3_address),                    //      .address
		.s0_write         (mw3_write),                      //      .write
		.s0_read          (mw3_read),                       //      .read
		.s0_byteenable    (mw3_byteenable),                 //      .byteenable
		.s0_debugaccess   (mw3_debugaccess),                //      .debugaccess
		.m0_waitrequest   (mm_bridge_9_m0_waitrequest),     //    m0.waitrequest
		.m0_readdata      (mm_bridge_9_m0_readdata),        //      .readdata
		.m0_readdatavalid (mm_bridge_9_m0_readdatavalid),   //      .readdatavalid
		.m0_burstcount    (mm_bridge_9_m0_burstcount),      //      .burstcount
		.m0_writedata     (mm_bridge_9_m0_writedata),       //      .writedata
		.m0_address       (mm_bridge_9_m0_address),         //      .address
		.m0_write         (mm_bridge_9_m0_write),           //      .write
		.m0_read          (mm_bridge_9_m0_read),            //      .read
		.m0_byteenable    (mm_bridge_9_m0_byteenable),      //      .byteenable
		.m0_debugaccess   (mm_bridge_9_m0_debugaccess)      //      .debugaccess
	);

	altera_avalon_mm_bridge #(
		.DATA_WIDTH        (128),
		.SYMBOL_WIDTH      (8),
		.ADDRESS_WIDTH     (26),
		.BURSTCOUNT_WIDTH  (6),
		.PIPELINE_COMMAND  (1),
		.PIPELINE_RESPONSE (1)
	) mm_bridge_10 (
		.clk              (hps_clk_clk),                        //   clk.clk
		.reset            (rst_controller_001_reset_out_reset), // reset.reset
		.s0_waitrequest   (hps_waitrequest),                    //    s0.waitrequest
		.s0_readdata      (hps_readdata),                       //      .readdata
		.s0_readdatavalid (hps_readdatavalid),                  //      .readdatavalid
		.s0_burstcount    (hps_burstcount),                     //      .burstcount
		.s0_writedata     (hps_writedata),                      //      .writedata
		.s0_address       (hps_address),                        //      .address
		.s0_write         (hps_write),                          //      .write
		.s0_read          (hps_read),                           //      .read
		.s0_byteenable    (hps_byteenable),                     //      .byteenable
		.s0_debugaccess   (hps_debugaccess),                    //      .debugaccess
		.m0_waitrequest   (mm_bridge_10_m0_waitrequest),        //    m0.waitrequest
		.m0_readdata      (mm_bridge_10_m0_readdata),           //      .readdata
		.m0_readdatavalid (mm_bridge_10_m0_readdatavalid),      //      .readdatavalid
		.m0_burstcount    (mm_bridge_10_m0_burstcount),         //      .burstcount
		.m0_writedata     (mm_bridge_10_m0_writedata),          //      .writedata
		.m0_address       (mm_bridge_10_m0_address),            //      .address
		.m0_write         (mm_bridge_10_m0_write),              //      .write
		.m0_read          (mm_bridge_10_m0_read),               //      .read
		.m0_byteenable    (mm_bridge_10_m0_byteenable),         //      .byteenable
		.m0_debugaccess   (mm_bridge_10_m0_debugaccess)         //      .debugaccess
	);

	altera_avalon_mm_bridge #(
		.DATA_WIDTH        (128),
		.SYMBOL_WIDTH      (8),
		.ADDRESS_WIDTH     (26),
		.BURSTCOUNT_WIDTH  (6),
		.PIPELINE_COMMAND  (1),
		.PIPELINE_RESPONSE (1)
	) mm_bridge_11 (
		.clk              (afi_clk_clk),                    //   clk.clk
		.reset            (rst_controller_reset_out_reset), // reset.reset
		.s0_waitrequest   (mwa_waitrequest),                //    s0.waitrequest
		.s0_readdata      (mwa_readdata),                   //      .readdata
		.s0_readdatavalid (mwa_readdatavalid),              //      .readdatavalid
		.s0_burstcount    (mwa_burstcount),                 //      .burstcount
		.s0_writedata     (mwa_writedata),                  //      .writedata
		.s0_address       (mwa_address),                    //      .address
		.s0_write         (mwa_write),                      //      .write
		.s0_read          (mwa_read),                       //      .read
		.s0_byteenable    (mwa_byteenable),                 //      .byteenable
		.s0_debugaccess   (mwa_debugaccess),                //      .debugaccess
		.m0_waitrequest   (mm_bridge_11_m0_waitrequest),    //    m0.waitrequest
		.m0_readdata      (mm_bridge_11_m0_readdata),       //      .readdata
		.m0_readdatavalid (mm_bridge_11_m0_readdatavalid),  //      .readdatavalid
		.m0_burstcount    (mm_bridge_11_m0_burstcount),     //      .burstcount
		.m0_writedata     (mm_bridge_11_m0_writedata),      //      .writedata
		.m0_address       (mm_bridge_11_m0_address),        //      .address
		.m0_write         (mm_bridge_11_m0_write),          //      .write
		.m0_read          (mm_bridge_11_m0_read),           //      .read
		.m0_byteenable    (mm_bridge_11_m0_byteenable),     //      .byteenable
		.m0_debugaccess   (mm_bridge_11_m0_debugaccess)     //      .debugaccess
	);

	fpga_mem_mm_interconnect_0 mm_interconnect_0 (
		.clock_bridge_1_out_clk_clk                                      (hps_clk_clk),                                                   //                                    clock_bridge_1_out_clk.clk
		.mem_if_ddr3_emif_0_afi_half_clk_clk                             (afi_clk_clk),                                                   //                           mem_if_ddr3_emif_0_afi_half_clk.clk
		.mem_if_ddr3_emif_0_mp_cmd_reset_n_0_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                                // mem_if_ddr3_emif_0_mp_cmd_reset_n_0_reset_bridge_in_reset.reset
		.mm_bridge_10_reset_reset_bridge_in_reset_reset                  (rst_controller_001_reset_out_reset),                            //                  mm_bridge_10_reset_reset_bridge_in_reset.reset
		.mm_bridge_11_reset_reset_bridge_in_reset_reset                  (rst_controller_reset_out_reset),                                //                  mm_bridge_11_reset_reset_bridge_in_reset.reset
		.mm_bridge_0_m0_address                                          (mm_bridge_0_m0_address),                                        //                                            mm_bridge_0_m0.address
		.mm_bridge_0_m0_waitrequest                                      (mm_bridge_0_m0_waitrequest),                                    //                                                          .waitrequest
		.mm_bridge_0_m0_burstcount                                       (mm_bridge_0_m0_burstcount),                                     //                                                          .burstcount
		.mm_bridge_0_m0_byteenable                                       (mm_bridge_0_m0_byteenable),                                     //                                                          .byteenable
		.mm_bridge_0_m0_read                                             (mm_bridge_0_m0_read),                                           //                                                          .read
		.mm_bridge_0_m0_readdata                                         (mm_bridge_0_m0_readdata),                                       //                                                          .readdata
		.mm_bridge_0_m0_readdatavalid                                    (mm_bridge_0_m0_readdatavalid),                                  //                                                          .readdatavalid
		.mm_bridge_0_m0_write                                            (mm_bridge_0_m0_write),                                          //                                                          .write
		.mm_bridge_0_m0_writedata                                        (mm_bridge_0_m0_writedata),                                      //                                                          .writedata
		.mm_bridge_0_m0_debugaccess                                      (mm_bridge_0_m0_debugaccess),                                    //                                                          .debugaccess
		.mm_bridge_1_m0_address                                          (mm_bridge_1_m0_address),                                        //                                            mm_bridge_1_m0.address
		.mm_bridge_1_m0_waitrequest                                      (mm_bridge_1_m0_waitrequest),                                    //                                                          .waitrequest
		.mm_bridge_1_m0_burstcount                                       (mm_bridge_1_m0_burstcount),                                     //                                                          .burstcount
		.mm_bridge_1_m0_byteenable                                       (mm_bridge_1_m0_byteenable),                                     //                                                          .byteenable
		.mm_bridge_1_m0_read                                             (mm_bridge_1_m0_read),                                           //                                                          .read
		.mm_bridge_1_m0_readdata                                         (mm_bridge_1_m0_readdata),                                       //                                                          .readdata
		.mm_bridge_1_m0_readdatavalid                                    (mm_bridge_1_m0_readdatavalid),                                  //                                                          .readdatavalid
		.mm_bridge_1_m0_write                                            (mm_bridge_1_m0_write),                                          //                                                          .write
		.mm_bridge_1_m0_writedata                                        (mm_bridge_1_m0_writedata),                                      //                                                          .writedata
		.mm_bridge_1_m0_debugaccess                                      (mm_bridge_1_m0_debugaccess),                                    //                                                          .debugaccess
		.mm_bridge_10_m0_address                                         (mm_bridge_10_m0_address),                                       //                                           mm_bridge_10_m0.address
		.mm_bridge_10_m0_waitrequest                                     (mm_bridge_10_m0_waitrequest),                                   //                                                          .waitrequest
		.mm_bridge_10_m0_burstcount                                      (mm_bridge_10_m0_burstcount),                                    //                                                          .burstcount
		.mm_bridge_10_m0_byteenable                                      (mm_bridge_10_m0_byteenable),                                    //                                                          .byteenable
		.mm_bridge_10_m0_read                                            (mm_bridge_10_m0_read),                                          //                                                          .read
		.mm_bridge_10_m0_readdata                                        (mm_bridge_10_m0_readdata),                                      //                                                          .readdata
		.mm_bridge_10_m0_readdatavalid                                   (mm_bridge_10_m0_readdatavalid),                                 //                                                          .readdatavalid
		.mm_bridge_10_m0_write                                           (mm_bridge_10_m0_write),                                         //                                                          .write
		.mm_bridge_10_m0_writedata                                       (mm_bridge_10_m0_writedata),                                     //                                                          .writedata
		.mm_bridge_10_m0_debugaccess                                     (mm_bridge_10_m0_debugaccess),                                   //                                                          .debugaccess
		.mm_bridge_11_m0_address                                         (mm_bridge_11_m0_address),                                       //                                           mm_bridge_11_m0.address
		.mm_bridge_11_m0_waitrequest                                     (mm_bridge_11_m0_waitrequest),                                   //                                                          .waitrequest
		.mm_bridge_11_m0_burstcount                                      (mm_bridge_11_m0_burstcount),                                    //                                                          .burstcount
		.mm_bridge_11_m0_byteenable                                      (mm_bridge_11_m0_byteenable),                                    //                                                          .byteenable
		.mm_bridge_11_m0_read                                            (mm_bridge_11_m0_read),                                          //                                                          .read
		.mm_bridge_11_m0_readdata                                        (mm_bridge_11_m0_readdata),                                      //                                                          .readdata
		.mm_bridge_11_m0_readdatavalid                                   (mm_bridge_11_m0_readdatavalid),                                 //                                                          .readdatavalid
		.mm_bridge_11_m0_write                                           (mm_bridge_11_m0_write),                                         //                                                          .write
		.mm_bridge_11_m0_writedata                                       (mm_bridge_11_m0_writedata),                                     //                                                          .writedata
		.mm_bridge_11_m0_debugaccess                                     (mm_bridge_11_m0_debugaccess),                                   //                                                          .debugaccess
		.mm_bridge_2_m0_address                                          (mm_bridge_2_m0_address),                                        //                                            mm_bridge_2_m0.address
		.mm_bridge_2_m0_waitrequest                                      (mm_bridge_2_m0_waitrequest),                                    //                                                          .waitrequest
		.mm_bridge_2_m0_burstcount                                       (mm_bridge_2_m0_burstcount),                                     //                                                          .burstcount
		.mm_bridge_2_m0_byteenable                                       (mm_bridge_2_m0_byteenable),                                     //                                                          .byteenable
		.mm_bridge_2_m0_read                                             (mm_bridge_2_m0_read),                                           //                                                          .read
		.mm_bridge_2_m0_readdata                                         (mm_bridge_2_m0_readdata),                                       //                                                          .readdata
		.mm_bridge_2_m0_readdatavalid                                    (mm_bridge_2_m0_readdatavalid),                                  //                                                          .readdatavalid
		.mm_bridge_2_m0_write                                            (mm_bridge_2_m0_write),                                          //                                                          .write
		.mm_bridge_2_m0_writedata                                        (mm_bridge_2_m0_writedata),                                      //                                                          .writedata
		.mm_bridge_2_m0_debugaccess                                      (mm_bridge_2_m0_debugaccess),                                    //                                                          .debugaccess
		.mm_bridge_3_m0_address                                          (mm_bridge_3_m0_address),                                        //                                            mm_bridge_3_m0.address
		.mm_bridge_3_m0_waitrequest                                      (mm_bridge_3_m0_waitrequest),                                    //                                                          .waitrequest
		.mm_bridge_3_m0_burstcount                                       (mm_bridge_3_m0_burstcount),                                     //                                                          .burstcount
		.mm_bridge_3_m0_byteenable                                       (mm_bridge_3_m0_byteenable),                                     //                                                          .byteenable
		.mm_bridge_3_m0_read                                             (mm_bridge_3_m0_read),                                           //                                                          .read
		.mm_bridge_3_m0_readdata                                         (mm_bridge_3_m0_readdata),                                       //                                                          .readdata
		.mm_bridge_3_m0_readdatavalid                                    (mm_bridge_3_m0_readdatavalid),                                  //                                                          .readdatavalid
		.mm_bridge_3_m0_write                                            (mm_bridge_3_m0_write),                                          //                                                          .write
		.mm_bridge_3_m0_writedata                                        (mm_bridge_3_m0_writedata),                                      //                                                          .writedata
		.mm_bridge_3_m0_debugaccess                                      (mm_bridge_3_m0_debugaccess),                                    //                                                          .debugaccess
		.mm_bridge_4_m0_address                                          (mm_bridge_4_m0_address),                                        //                                            mm_bridge_4_m0.address
		.mm_bridge_4_m0_waitrequest                                      (mm_bridge_4_m0_waitrequest),                                    //                                                          .waitrequest
		.mm_bridge_4_m0_burstcount                                       (mm_bridge_4_m0_burstcount),                                     //                                                          .burstcount
		.mm_bridge_4_m0_byteenable                                       (mm_bridge_4_m0_byteenable),                                     //                                                          .byteenable
		.mm_bridge_4_m0_read                                             (mm_bridge_4_m0_read),                                           //                                                          .read
		.mm_bridge_4_m0_readdata                                         (mm_bridge_4_m0_readdata),                                       //                                                          .readdata
		.mm_bridge_4_m0_readdatavalid                                    (mm_bridge_4_m0_readdatavalid),                                  //                                                          .readdatavalid
		.mm_bridge_4_m0_write                                            (mm_bridge_4_m0_write),                                          //                                                          .write
		.mm_bridge_4_m0_writedata                                        (mm_bridge_4_m0_writedata),                                      //                                                          .writedata
		.mm_bridge_4_m0_debugaccess                                      (mm_bridge_4_m0_debugaccess),                                    //                                                          .debugaccess
		.mm_bridge_5_m0_address                                          (mm_bridge_5_m0_address),                                        //                                            mm_bridge_5_m0.address
		.mm_bridge_5_m0_waitrequest                                      (mm_bridge_5_m0_waitrequest),                                    //                                                          .waitrequest
		.mm_bridge_5_m0_burstcount                                       (mm_bridge_5_m0_burstcount),                                     //                                                          .burstcount
		.mm_bridge_5_m0_byteenable                                       (mm_bridge_5_m0_byteenable),                                     //                                                          .byteenable
		.mm_bridge_5_m0_read                                             (mm_bridge_5_m0_read),                                           //                                                          .read
		.mm_bridge_5_m0_readdata                                         (mm_bridge_5_m0_readdata),                                       //                                                          .readdata
		.mm_bridge_5_m0_readdatavalid                                    (mm_bridge_5_m0_readdatavalid),                                  //                                                          .readdatavalid
		.mm_bridge_5_m0_write                                            (mm_bridge_5_m0_write),                                          //                                                          .write
		.mm_bridge_5_m0_writedata                                        (mm_bridge_5_m0_writedata),                                      //                                                          .writedata
		.mm_bridge_5_m0_debugaccess                                      (mm_bridge_5_m0_debugaccess),                                    //                                                          .debugaccess
		.mm_bridge_6_m0_address                                          (mm_bridge_6_m0_address),                                        //                                            mm_bridge_6_m0.address
		.mm_bridge_6_m0_waitrequest                                      (mm_bridge_6_m0_waitrequest),                                    //                                                          .waitrequest
		.mm_bridge_6_m0_burstcount                                       (mm_bridge_6_m0_burstcount),                                     //                                                          .burstcount
		.mm_bridge_6_m0_byteenable                                       (mm_bridge_6_m0_byteenable),                                     //                                                          .byteenable
		.mm_bridge_6_m0_read                                             (mm_bridge_6_m0_read),                                           //                                                          .read
		.mm_bridge_6_m0_readdata                                         (mm_bridge_6_m0_readdata),                                       //                                                          .readdata
		.mm_bridge_6_m0_readdatavalid                                    (mm_bridge_6_m0_readdatavalid),                                  //                                                          .readdatavalid
		.mm_bridge_6_m0_write                                            (mm_bridge_6_m0_write),                                          //                                                          .write
		.mm_bridge_6_m0_writedata                                        (mm_bridge_6_m0_writedata),                                      //                                                          .writedata
		.mm_bridge_6_m0_debugaccess                                      (mm_bridge_6_m0_debugaccess),                                    //                                                          .debugaccess
		.mm_bridge_7_m0_address                                          (mm_bridge_7_m0_address),                                        //                                            mm_bridge_7_m0.address
		.mm_bridge_7_m0_waitrequest                                      (mm_bridge_7_m0_waitrequest),                                    //                                                          .waitrequest
		.mm_bridge_7_m0_burstcount                                       (mm_bridge_7_m0_burstcount),                                     //                                                          .burstcount
		.mm_bridge_7_m0_byteenable                                       (mm_bridge_7_m0_byteenable),                                     //                                                          .byteenable
		.mm_bridge_7_m0_read                                             (mm_bridge_7_m0_read),                                           //                                                          .read
		.mm_bridge_7_m0_readdata                                         (mm_bridge_7_m0_readdata),                                       //                                                          .readdata
		.mm_bridge_7_m0_readdatavalid                                    (mm_bridge_7_m0_readdatavalid),                                  //                                                          .readdatavalid
		.mm_bridge_7_m0_write                                            (mm_bridge_7_m0_write),                                          //                                                          .write
		.mm_bridge_7_m0_writedata                                        (mm_bridge_7_m0_writedata),                                      //                                                          .writedata
		.mm_bridge_7_m0_debugaccess                                      (mm_bridge_7_m0_debugaccess),                                    //                                                          .debugaccess
		.mm_bridge_8_m0_address                                          (mm_bridge_8_m0_address),                                        //                                            mm_bridge_8_m0.address
		.mm_bridge_8_m0_waitrequest                                      (mm_bridge_8_m0_waitrequest),                                    //                                                          .waitrequest
		.mm_bridge_8_m0_burstcount                                       (mm_bridge_8_m0_burstcount),                                     //                                                          .burstcount
		.mm_bridge_8_m0_byteenable                                       (mm_bridge_8_m0_byteenable),                                     //                                                          .byteenable
		.mm_bridge_8_m0_read                                             (mm_bridge_8_m0_read),                                           //                                                          .read
		.mm_bridge_8_m0_readdata                                         (mm_bridge_8_m0_readdata),                                       //                                                          .readdata
		.mm_bridge_8_m0_readdatavalid                                    (mm_bridge_8_m0_readdatavalid),                                  //                                                          .readdatavalid
		.mm_bridge_8_m0_write                                            (mm_bridge_8_m0_write),                                          //                                                          .write
		.mm_bridge_8_m0_writedata                                        (mm_bridge_8_m0_writedata),                                      //                                                          .writedata
		.mm_bridge_8_m0_debugaccess                                      (mm_bridge_8_m0_debugaccess),                                    //                                                          .debugaccess
		.mm_bridge_9_m0_address                                          (mm_bridge_9_m0_address),                                        //                                            mm_bridge_9_m0.address
		.mm_bridge_9_m0_waitrequest                                      (mm_bridge_9_m0_waitrequest),                                    //                                                          .waitrequest
		.mm_bridge_9_m0_burstcount                                       (mm_bridge_9_m0_burstcount),                                     //                                                          .burstcount
		.mm_bridge_9_m0_byteenable                                       (mm_bridge_9_m0_byteenable),                                     //                                                          .byteenable
		.mm_bridge_9_m0_read                                             (mm_bridge_9_m0_read),                                           //                                                          .read
		.mm_bridge_9_m0_readdata                                         (mm_bridge_9_m0_readdata),                                       //                                                          .readdata
		.mm_bridge_9_m0_readdatavalid                                    (mm_bridge_9_m0_readdatavalid),                                  //                                                          .readdatavalid
		.mm_bridge_9_m0_write                                            (mm_bridge_9_m0_write),                                          //                                                          .write
		.mm_bridge_9_m0_writedata                                        (mm_bridge_9_m0_writedata),                                      //                                                          .writedata
		.mm_bridge_9_m0_debugaccess                                      (mm_bridge_9_m0_debugaccess),                                    //                                                          .debugaccess
		.mem_if_ddr3_emif_0_avl_0_address                                (mm_interconnect_0_mem_if_ddr3_emif_0_avl_0_address),            //                                  mem_if_ddr3_emif_0_avl_0.address
		.mem_if_ddr3_emif_0_avl_0_write                                  (mm_interconnect_0_mem_if_ddr3_emif_0_avl_0_write),              //                                                          .write
		.mem_if_ddr3_emif_0_avl_0_read                                   (mm_interconnect_0_mem_if_ddr3_emif_0_avl_0_read),               //                                                          .read
		.mem_if_ddr3_emif_0_avl_0_readdata                               (mm_interconnect_0_mem_if_ddr3_emif_0_avl_0_readdata),           //                                                          .readdata
		.mem_if_ddr3_emif_0_avl_0_writedata                              (mm_interconnect_0_mem_if_ddr3_emif_0_avl_0_writedata),          //                                                          .writedata
		.mem_if_ddr3_emif_0_avl_0_beginbursttransfer                     (mm_interconnect_0_mem_if_ddr3_emif_0_avl_0_beginbursttransfer), //                                                          .beginbursttransfer
		.mem_if_ddr3_emif_0_avl_0_burstcount                             (mm_interconnect_0_mem_if_ddr3_emif_0_avl_0_burstcount),         //                                                          .burstcount
		.mem_if_ddr3_emif_0_avl_0_byteenable                             (mm_interconnect_0_mem_if_ddr3_emif_0_avl_0_byteenable),         //                                                          .byteenable
		.mem_if_ddr3_emif_0_avl_0_readdatavalid                          (mm_interconnect_0_mem_if_ddr3_emif_0_avl_0_readdatavalid),      //                                                          .readdatavalid
		.mem_if_ddr3_emif_0_avl_0_waitrequest                            (~mm_interconnect_0_mem_if_ddr3_emif_0_avl_0_waitrequest)        //                                                          .waitrequest
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                 // reset_in0.reset
		.clk            (afi_clk_clk),                    //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (hps_clk_clk),                        //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
