// soc_system_tb.v

// Generated using ACDS version 13.1 162 at 2015.06.22.13:03:10

`timescale 1 ps / 1 ps
module soc_system_tb (
	);

	wire          soc_system_inst_clk_bfm_clk_clk;                                   // soc_system_inst_clk_bfm:clk -> [soc_system_inst:clk_clk, soc_system_inst_hps_0_f2h_cold_reset_req_bfm:clk, soc_system_inst_hps_0_f2h_debug_reset_req_bfm:clk, soc_system_inst_hps_0_f2h_warm_reset_req_bfm:clk, soc_system_inst_reg_avl_bfm:clk, soc_system_inst_reset_bfm:clk]
	wire          soc_system_inst_afi_clk_bfm_clk_clk;                               // soc_system_inst_afi_clk_bfm:clk -> [rst_controller:clk, soc_system_inst:afi_clk_clk, soc_system_inst_h2f_0_bfm:clk]
	wire          soc_system_inst_reset_bfm_reset_reset;                             // soc_system_inst_reset_bfm:reset -> [rst_controller:reset_in0, soc_system_inst:reset_reset_n, soc_system_inst_reg_avl_bfm:reset]
	wire          soc_system_inst_hps_0_f2h_warm_reset_req_bfm_reset_reset;          // soc_system_inst_hps_0_f2h_warm_reset_req_bfm:reset -> soc_system_inst:hps_0_f2h_warm_reset_req_reset_n
	wire          soc_system_inst_hps_0_f2h_debug_reset_req_bfm_reset_reset;         // soc_system_inst_hps_0_f2h_debug_reset_req_bfm:reset -> soc_system_inst:hps_0_f2h_debug_reset_req_reset_n
	wire          soc_system_inst_hps_0_f2h_cold_reset_req_bfm_reset_reset;          // soc_system_inst_hps_0_f2h_cold_reset_req_bfm:reset -> soc_system_inst:hps_0_f2h_cold_reset_req_reset_n
	wire          soc_system_inst_memory_mem_odt;                                    // soc_system_inst:memory_mem_odt -> soc_system_inst_memory_bfm:sig_mem_odt
	wire          soc_system_inst_memory_mem_cs_n;                                   // soc_system_inst:memory_mem_cs_n -> soc_system_inst_memory_bfm:sig_mem_cs_n
	wire   [14:0] soc_system_inst_memory_mem_a;                                      // soc_system_inst:memory_mem_a -> soc_system_inst_memory_bfm:sig_mem_a
	wire    [0:0] soc_system_inst_memory_bfm_conduit_oct_rzqin;                      // soc_system_inst_memory_bfm:sig_oct_rzqin -> soc_system_inst:memory_oct_rzqin
	wire          soc_system_inst_memory_mem_ck_n;                                   // soc_system_inst:memory_mem_ck_n -> soc_system_inst_memory_bfm:sig_mem_ck_n
	wire          soc_system_inst_memory_mem_ras_n;                                  // soc_system_inst:memory_mem_ras_n -> soc_system_inst_memory_bfm:sig_mem_ras_n
	wire          soc_system_inst_memory_mem_cke;                                    // soc_system_inst:memory_mem_cke -> soc_system_inst_memory_bfm:sig_mem_cke
	wire    [3:0] soc_system_inst_memory_mem_dqs;                                    // [] -> [soc_system_inst:memory_mem_dqs, soc_system_inst_memory_bfm:sig_mem_dqs]
	wire          soc_system_inst_memory_mem_we_n;                                   // soc_system_inst:memory_mem_we_n -> soc_system_inst_memory_bfm:sig_mem_we_n
	wire    [2:0] soc_system_inst_memory_mem_ba;                                     // soc_system_inst:memory_mem_ba -> soc_system_inst_memory_bfm:sig_mem_ba
	wire   [31:0] soc_system_inst_memory_mem_dq;                                     // [] -> [soc_system_inst:memory_mem_dq, soc_system_inst_memory_bfm:sig_mem_dq]
	wire          soc_system_inst_memory_mem_ck;                                     // soc_system_inst:memory_mem_ck -> soc_system_inst_memory_bfm:sig_mem_ck
	wire          soc_system_inst_memory_mem_reset_n;                                // soc_system_inst:memory_mem_reset_n -> soc_system_inst_memory_bfm:sig_mem_reset_n
	wire    [3:0] soc_system_inst_memory_mem_dm;                                     // soc_system_inst:memory_mem_dm -> soc_system_inst_memory_bfm:sig_mem_dm
	wire          soc_system_inst_memory_mem_cas_n;                                  // soc_system_inst:memory_mem_cas_n -> soc_system_inst_memory_bfm:sig_mem_cas_n
	wire    [3:0] soc_system_inst_memory_mem_dqs_n;                                  // [] -> [soc_system_inst:memory_mem_dqs_n, soc_system_inst_memory_bfm:sig_mem_dqs_n]
	wire          soc_system_inst_hps_0_hps_io_hps_io_gpio_inst_gpio35;              // [] -> [soc_system_inst:hps_0_hps_io_hps_io_gpio_inst_GPIO35, soc_system_inst_hps_0_hps_io_bfm:sig_hps_io_gpio_inst_GPIO35]
	wire          soc_system_inst_hps_0_hps_io_hps_io_emac1_inst_tx_ctl;             // soc_system_inst:hps_0_hps_io_hps_io_emac1_inst_TX_CTL -> soc_system_inst_hps_0_hps_io_bfm:sig_hps_io_emac1_inst_TX_CTL
	wire          soc_system_inst_hps_0_hps_io_hps_io_emac1_inst_mdio;               // [] -> [soc_system_inst:hps_0_hps_io_hps_io_emac1_inst_MDIO, soc_system_inst_hps_0_hps_io_bfm:sig_hps_io_emac1_inst_MDIO]
	wire          soc_system_inst_hps_0_hps_io_hps_io_spim0_inst_mosi;               // soc_system_inst:hps_0_hps_io_hps_io_spim0_inst_MOSI -> soc_system_inst_hps_0_hps_io_bfm:sig_hps_io_spim0_inst_MOSI
	wire          soc_system_inst_hps_0_hps_io_hps_io_gpio_inst_gpio62;              // [] -> [soc_system_inst:hps_0_hps_io_hps_io_gpio_inst_GPIO62, soc_system_inst_hps_0_hps_io_bfm:sig_hps_io_gpio_inst_GPIO62]
	wire          soc_system_inst_hps_0_hps_io_hps_io_gpio_inst_gpio61;              // [] -> [soc_system_inst:hps_0_hps_io_hps_io_gpio_inst_GPIO61, soc_system_inst_hps_0_hps_io_bfm:sig_hps_io_gpio_inst_GPIO61]
	wire          soc_system_inst_hps_0_hps_io_hps_io_usb1_inst_d5;                  // [] -> [soc_system_inst:hps_0_hps_io_hps_io_usb1_inst_D5, soc_system_inst_hps_0_hps_io_bfm:sig_hps_io_usb1_inst_D5]
	wire    [0:0] soc_system_inst_hps_0_hps_io_bfm_conduit_hps_io_usb1_inst_clk;     // soc_system_inst_hps_0_hps_io_bfm:sig_hps_io_usb1_inst_CLK -> soc_system_inst:hps_0_hps_io_hps_io_usb1_inst_CLK
	wire    [0:0] soc_system_inst_hps_0_hps_io_bfm_conduit_hps_io_spim1_inst_miso;   // soc_system_inst_hps_0_hps_io_bfm:sig_hps_io_spim1_inst_MISO -> soc_system_inst:hps_0_hps_io_hps_io_spim1_inst_MISO
	wire          soc_system_inst_hps_0_hps_io_hps_io_usb1_inst_d4;                  // [] -> [soc_system_inst:hps_0_hps_io_hps_io_usb1_inst_D4, soc_system_inst_hps_0_hps_io_bfm:sig_hps_io_usb1_inst_D4]
	wire          soc_system_inst_hps_0_hps_io_hps_io_usb1_inst_d7;                  // [] -> [soc_system_inst:hps_0_hps_io_hps_io_usb1_inst_D7, soc_system_inst_hps_0_hps_io_bfm:sig_hps_io_usb1_inst_D7]
	wire          soc_system_inst_hps_0_hps_io_hps_io_usb1_inst_d6;                  // [] -> [soc_system_inst:hps_0_hps_io_hps_io_usb1_inst_D6, soc_system_inst_hps_0_hps_io_bfm:sig_hps_io_usb1_inst_D6]
	wire          soc_system_inst_hps_0_hps_io_hps_io_usb1_inst_d1;                  // [] -> [soc_system_inst:hps_0_hps_io_hps_io_usb1_inst_D1, soc_system_inst_hps_0_hps_io_bfm:sig_hps_io_usb1_inst_D1]
	wire          soc_system_inst_hps_0_hps_io_hps_io_usb1_inst_d0;                  // [] -> [soc_system_inst:hps_0_hps_io_hps_io_usb1_inst_D0, soc_system_inst_hps_0_hps_io_bfm:sig_hps_io_usb1_inst_D0]
	wire          soc_system_inst_hps_0_hps_io_hps_io_usb1_inst_d3;                  // [] -> [soc_system_inst:hps_0_hps_io_hps_io_usb1_inst_D3, soc_system_inst_hps_0_hps_io_bfm:sig_hps_io_usb1_inst_D3]
	wire    [0:0] soc_system_inst_hps_0_hps_io_bfm_conduit_hps_io_emac1_inst_rx_clk; // soc_system_inst_hps_0_hps_io_bfm:sig_hps_io_emac1_inst_RX_CLK -> soc_system_inst:hps_0_hps_io_hps_io_emac1_inst_RX_CLK
	wire          soc_system_inst_hps_0_hps_io_hps_io_usb1_inst_d2;                  // [] -> [soc_system_inst:hps_0_hps_io_hps_io_usb1_inst_D2, soc_system_inst_hps_0_hps_io_bfm:sig_hps_io_usb1_inst_D2]
	wire    [0:0] soc_system_inst_hps_0_hps_io_bfm_conduit_hps_io_uart0_inst_rx;     // soc_system_inst_hps_0_hps_io_bfm:sig_hps_io_uart0_inst_RX -> soc_system_inst:hps_0_hps_io_hps_io_uart0_inst_RX
	wire          soc_system_inst_hps_0_hps_io_hps_io_spim1_inst_ss0;                // soc_system_inst:hps_0_hps_io_hps_io_spim1_inst_SS0 -> soc_system_inst_hps_0_hps_io_bfm:sig_hps_io_spim1_inst_SS0
	wire          soc_system_inst_hps_0_hps_io_hps_io_spim0_inst_ss0;                // soc_system_inst:hps_0_hps_io_hps_io_spim0_inst_SS0 -> soc_system_inst_hps_0_hps_io_bfm:sig_hps_io_spim0_inst_SS0
	wire    [0:0] soc_system_inst_hps_0_hps_io_bfm_conduit_hps_io_emac1_inst_rxd3;   // soc_system_inst_hps_0_hps_io_bfm:sig_hps_io_emac1_inst_RXD3 -> soc_system_inst:hps_0_hps_io_hps_io_emac1_inst_RXD3
	wire    [0:0] soc_system_inst_hps_0_hps_io_bfm_conduit_hps_io_emac1_inst_rxd2;   // soc_system_inst_hps_0_hps_io_bfm:sig_hps_io_emac1_inst_RXD2 -> soc_system_inst:hps_0_hps_io_hps_io_emac1_inst_RXD2
	wire          soc_system_inst_hps_0_hps_io_hps_io_i2c1_inst_scl;                 // [] -> [soc_system_inst:hps_0_hps_io_hps_io_i2c1_inst_SCL, soc_system_inst_hps_0_hps_io_bfm:sig_hps_io_i2c1_inst_SCL]
	wire    [0:0] soc_system_inst_hps_0_hps_io_bfm_conduit_hps_io_emac1_inst_rx_ctl; // soc_system_inst_hps_0_hps_io_bfm:sig_hps_io_emac1_inst_RX_CTL -> soc_system_inst:hps_0_hps_io_hps_io_emac1_inst_RX_CTL
	wire          soc_system_inst_hps_0_hps_io_hps_io_usb1_inst_stp;                 // soc_system_inst:hps_0_hps_io_hps_io_usb1_inst_STP -> soc_system_inst_hps_0_hps_io_bfm:sig_hps_io_usb1_inst_STP
	wire          soc_system_inst_hps_0_hps_io_hps_io_sdio_inst_clk;                 // soc_system_inst:hps_0_hps_io_hps_io_sdio_inst_CLK -> soc_system_inst_hps_0_hps_io_bfm:sig_hps_io_sdio_inst_CLK
	wire          soc_system_inst_hps_0_hps_io_hps_io_sdio_inst_d1;                  // [] -> [soc_system_inst:hps_0_hps_io_hps_io_sdio_inst_D1, soc_system_inst_hps_0_hps_io_bfm:sig_hps_io_sdio_inst_D1]
	wire          soc_system_inst_hps_0_hps_io_hps_io_gpio_inst_gpio53;              // [] -> [soc_system_inst:hps_0_hps_io_hps_io_gpio_inst_GPIO53, soc_system_inst_hps_0_hps_io_bfm:sig_hps_io_gpio_inst_GPIO53]
	wire          soc_system_inst_hps_0_hps_io_hps_io_sdio_inst_d0;                  // [] -> [soc_system_inst:hps_0_hps_io_hps_io_sdio_inst_D0, soc_system_inst_hps_0_hps_io_bfm:sig_hps_io_sdio_inst_D0]
	wire          soc_system_inst_hps_0_hps_io_hps_io_gpio_inst_gpio54;              // [] -> [soc_system_inst:hps_0_hps_io_hps_io_gpio_inst_GPIO54, soc_system_inst_hps_0_hps_io_bfm:sig_hps_io_gpio_inst_GPIO54]
	wire          soc_system_inst_hps_0_hps_io_hps_io_sdio_inst_d3;                  // [] -> [soc_system_inst:hps_0_hps_io_hps_io_sdio_inst_D3, soc_system_inst_hps_0_hps_io_bfm:sig_hps_io_sdio_inst_D3]
	wire          soc_system_inst_hps_0_hps_io_hps_io_gpio_inst_gpio55;              // [] -> [soc_system_inst:hps_0_hps_io_hps_io_gpio_inst_GPIO55, soc_system_inst_hps_0_hps_io_bfm:sig_hps_io_gpio_inst_GPIO55]
	wire          soc_system_inst_hps_0_hps_io_hps_io_sdio_inst_d2;                  // [] -> [soc_system_inst:hps_0_hps_io_hps_io_sdio_inst_D2, soc_system_inst_hps_0_hps_io_bfm:sig_hps_io_sdio_inst_D2]
	wire          soc_system_inst_hps_0_hps_io_hps_io_gpio_inst_gpio56;              // [] -> [soc_system_inst:hps_0_hps_io_hps_io_gpio_inst_GPIO56, soc_system_inst_hps_0_hps_io_bfm:sig_hps_io_gpio_inst_GPIO56]
	wire    [0:0] soc_system_inst_hps_0_hps_io_bfm_conduit_hps_io_spim0_inst_miso;   // soc_system_inst_hps_0_hps_io_bfm:sig_hps_io_spim0_inst_MISO -> soc_system_inst:hps_0_hps_io_hps_io_spim0_inst_MISO
	wire          soc_system_inst_hps_0_hps_io_hps_io_gpio_inst_gpio48;              // [] -> [soc_system_inst:hps_0_hps_io_hps_io_gpio_inst_GPIO48, soc_system_inst_hps_0_hps_io_bfm:sig_hps_io_gpio_inst_GPIO48]
	wire          soc_system_inst_hps_0_hps_io_hps_io_gpio_inst_gpio00;              // [] -> [soc_system_inst:hps_0_hps_io_hps_io_gpio_inst_GPIO00, soc_system_inst_hps_0_hps_io_bfm:sig_hps_io_gpio_inst_GPIO00]
	wire          soc_system_inst_hps_0_hps_io_hps_io_qspi_inst_io3;                 // [] -> [soc_system_inst:hps_0_hps_io_hps_io_qspi_inst_IO3, soc_system_inst_hps_0_hps_io_bfm:sig_hps_io_qspi_inst_IO3]
	wire          soc_system_inst_hps_0_hps_io_hps_io_emac1_inst_txd1;               // soc_system_inst:hps_0_hps_io_hps_io_emac1_inst_TXD1 -> soc_system_inst_hps_0_hps_io_bfm:sig_hps_io_emac1_inst_TXD1
	wire          soc_system_inst_hps_0_hps_io_hps_io_qspi_inst_io2;                 // [] -> [soc_system_inst:hps_0_hps_io_hps_io_qspi_inst_IO2, soc_system_inst_hps_0_hps_io_bfm:sig_hps_io_qspi_inst_IO2]
	wire          soc_system_inst_hps_0_hps_io_hps_io_emac1_inst_txd0;               // soc_system_inst:hps_0_hps_io_hps_io_emac1_inst_TXD0 -> soc_system_inst_hps_0_hps_io_bfm:sig_hps_io_emac1_inst_TXD0
	wire          soc_system_inst_hps_0_hps_io_hps_io_qspi_inst_io1;                 // [] -> [soc_system_inst:hps_0_hps_io_hps_io_qspi_inst_IO1, soc_system_inst_hps_0_hps_io_bfm:sig_hps_io_qspi_inst_IO1]
	wire          soc_system_inst_hps_0_hps_io_hps_io_emac1_inst_txd3;               // soc_system_inst:hps_0_hps_io_hps_io_emac1_inst_TXD3 -> soc_system_inst_hps_0_hps_io_bfm:sig_hps_io_emac1_inst_TXD3
	wire          soc_system_inst_hps_0_hps_io_hps_io_qspi_inst_io0;                 // [] -> [soc_system_inst:hps_0_hps_io_hps_io_qspi_inst_IO0, soc_system_inst_hps_0_hps_io_bfm:sig_hps_io_qspi_inst_IO0]
	wire          soc_system_inst_hps_0_hps_io_hps_io_emac1_inst_txd2;               // soc_system_inst:hps_0_hps_io_hps_io_emac1_inst_TXD2 -> soc_system_inst_hps_0_hps_io_bfm:sig_hps_io_emac1_inst_TXD2
	wire    [0:0] soc_system_inst_hps_0_hps_io_bfm_conduit_hps_io_usb1_inst_dir;     // soc_system_inst_hps_0_hps_io_bfm:sig_hps_io_usb1_inst_DIR -> soc_system_inst:hps_0_hps_io_hps_io_usb1_inst_DIR
	wire    [0:0] soc_system_inst_hps_0_hps_io_bfm_conduit_hps_io_emac1_inst_rxd0;   // soc_system_inst_hps_0_hps_io_bfm:sig_hps_io_emac1_inst_RXD0 -> soc_system_inst:hps_0_hps_io_hps_io_emac1_inst_RXD0
	wire          soc_system_inst_hps_0_hps_io_hps_io_spim1_inst_clk;                // soc_system_inst:hps_0_hps_io_hps_io_spim1_inst_CLK -> soc_system_inst_hps_0_hps_io_bfm:sig_hps_io_spim1_inst_CLK
	wire          soc_system_inst_hps_0_hps_io_hps_io_i2c1_inst_sda;                 // [] -> [soc_system_inst:hps_0_hps_io_hps_io_i2c1_inst_SDA, soc_system_inst_hps_0_hps_io_bfm:sig_hps_io_i2c1_inst_SDA]
	wire    [0:0] soc_system_inst_hps_0_hps_io_bfm_conduit_hps_io_emac1_inst_rxd1;   // soc_system_inst_hps_0_hps_io_bfm:sig_hps_io_emac1_inst_RXD1 -> soc_system_inst:hps_0_hps_io_hps_io_emac1_inst_RXD1
	wire          soc_system_inst_hps_0_hps_io_hps_io_spim0_inst_clk;                // soc_system_inst:hps_0_hps_io_hps_io_spim0_inst_CLK -> soc_system_inst_hps_0_hps_io_bfm:sig_hps_io_spim0_inst_CLK
	wire          soc_system_inst_hps_0_hps_io_hps_io_sdio_inst_cmd;                 // [] -> [soc_system_inst:hps_0_hps_io_hps_io_sdio_inst_CMD, soc_system_inst_hps_0_hps_io_bfm:sig_hps_io_sdio_inst_CMD]
	wire          soc_system_inst_hps_0_hps_io_hps_io_qspi_inst_clk;                 // soc_system_inst:hps_0_hps_io_hps_io_qspi_inst_CLK -> soc_system_inst_hps_0_hps_io_bfm:sig_hps_io_qspi_inst_CLK
	wire          soc_system_inst_hps_0_hps_io_hps_io_gpio_inst_gpio09;              // [] -> [soc_system_inst:hps_0_hps_io_hps_io_gpio_inst_GPIO09, soc_system_inst_hps_0_hps_io_bfm:sig_hps_io_gpio_inst_GPIO09]
	wire          soc_system_inst_hps_0_hps_io_hps_io_gpio_inst_gpio40;              // [] -> [soc_system_inst:hps_0_hps_io_hps_io_gpio_inst_GPIO40, soc_system_inst_hps_0_hps_io_bfm:sig_hps_io_gpio_inst_GPIO40]
	wire          soc_system_inst_hps_0_hps_io_hps_io_emac1_inst_mdc;                // soc_system_inst:hps_0_hps_io_hps_io_emac1_inst_MDC -> soc_system_inst_hps_0_hps_io_bfm:sig_hps_io_emac1_inst_MDC
	wire          soc_system_inst_hps_0_hps_io_hps_io_uart0_inst_tx;                 // soc_system_inst:hps_0_hps_io_hps_io_uart0_inst_TX -> soc_system_inst_hps_0_hps_io_bfm:sig_hps_io_uart0_inst_TX
	wire    [0:0] soc_system_inst_hps_0_hps_io_bfm_conduit_hps_io_usb1_inst_nxt;     // soc_system_inst_hps_0_hps_io_bfm:sig_hps_io_usb1_inst_NXT -> soc_system_inst:hps_0_hps_io_hps_io_usb1_inst_NXT
	wire          soc_system_inst_hps_0_hps_io_hps_io_spim1_inst_mosi;               // soc_system_inst:hps_0_hps_io_hps_io_spim1_inst_MOSI -> soc_system_inst_hps_0_hps_io_bfm:sig_hps_io_spim1_inst_MOSI
	wire          soc_system_inst_hps_0_hps_io_hps_io_emac1_inst_tx_clk;             // soc_system_inst:hps_0_hps_io_hps_io_emac1_inst_TX_CLK -> soc_system_inst_hps_0_hps_io_bfm:sig_hps_io_emac1_inst_TX_CLK
	wire          soc_system_inst_hps_0_hps_io_hps_io_qspi_inst_ss0;                 // soc_system_inst:hps_0_hps_io_hps_io_qspi_inst_SS0 -> soc_system_inst_hps_0_hps_io_bfm:sig_hps_io_qspi_inst_SS0
	wire   [27:0] soc_system_inst_hps_0_f2h_stm_hw_events_bfm_conduit_stm_hwevents;  // soc_system_inst_hps_0_f2h_stm_hw_events_bfm:sig_stm_hwevents -> soc_system_inst:hps_0_f2h_stm_hw_events_stm_hwevents
	wire    [0:0] soc_system_inst_reg_avl_burstcount;                                // soc_system_inst:reg_avl_burstcount -> soc_system_inst_reg_avl_bfm:avs_burstcount
	wire          soc_system_inst_reg_avl_waitrequest;                               // soc_system_inst_reg_avl_bfm:avs_waitrequest -> soc_system_inst:reg_avl_waitrequest
	wire    [9:0] soc_system_inst_reg_avl_address;                                   // soc_system_inst:reg_avl_address -> soc_system_inst_reg_avl_bfm:avs_address
	wire   [31:0] soc_system_inst_reg_avl_writedata;                                 // soc_system_inst:reg_avl_writedata -> soc_system_inst_reg_avl_bfm:avs_writedata
	wire          soc_system_inst_reg_avl_write;                                     // soc_system_inst:reg_avl_write -> soc_system_inst_reg_avl_bfm:avs_write
	wire          soc_system_inst_reg_avl_read;                                      // soc_system_inst:reg_avl_read -> soc_system_inst_reg_avl_bfm:avs_read
	wire   [31:0] soc_system_inst_reg_avl_readdata;                                  // soc_system_inst_reg_avl_bfm:avs_readdata -> soc_system_inst:reg_avl_readdata
	wire          soc_system_inst_reg_avl_debugaccess;                               // soc_system_inst:reg_avl_debugaccess -> soc_system_inst_reg_avl_bfm:avs_debugaccess
	wire    [3:0] soc_system_inst_reg_avl_byteenable;                                // soc_system_inst:reg_avl_byteenable -> soc_system_inst_reg_avl_bfm:avs_byteenable
	wire          soc_system_inst_reg_avl_readdatavalid;                             // soc_system_inst_reg_avl_bfm:avs_readdatavalid -> soc_system_inst:reg_avl_readdatavalid
	wire    [5:0] soc_system_inst_h2f_0_burstcount;                                  // soc_system_inst:h2f_0_burstcount -> soc_system_inst_h2f_0_bfm:avs_burstcount
	wire          soc_system_inst_h2f_0_waitrequest;                                 // soc_system_inst_h2f_0_bfm:avs_waitrequest -> soc_system_inst:h2f_0_waitrequest
	wire   [25:0] soc_system_inst_h2f_0_address;                                     // soc_system_inst:h2f_0_address -> soc_system_inst_h2f_0_bfm:avs_address
	wire  [127:0] soc_system_inst_h2f_0_writedata;                                   // soc_system_inst:h2f_0_writedata -> soc_system_inst_h2f_0_bfm:avs_writedata
	wire          soc_system_inst_h2f_0_write;                                       // soc_system_inst:h2f_0_write -> soc_system_inst_h2f_0_bfm:avs_write
	wire          soc_system_inst_h2f_0_read;                                        // soc_system_inst:h2f_0_read -> soc_system_inst_h2f_0_bfm:avs_read
	wire  [127:0] soc_system_inst_h2f_0_readdata;                                    // soc_system_inst_h2f_0_bfm:avs_readdata -> soc_system_inst:h2f_0_readdata
	wire          soc_system_inst_h2f_0_debugaccess;                                 // soc_system_inst:h2f_0_debugaccess -> soc_system_inst_h2f_0_bfm:avs_debugaccess
	wire   [15:0] soc_system_inst_h2f_0_byteenable;                                  // soc_system_inst:h2f_0_byteenable -> soc_system_inst_h2f_0_bfm:avs_byteenable
	wire          soc_system_inst_h2f_0_readdatavalid;                               // soc_system_inst_h2f_0_bfm:avs_readdatavalid -> soc_system_inst:h2f_0_readdatavalid
	wire          rst_controller_reset_out_reset;                                    // rst_controller:reset_out -> soc_system_inst_h2f_0_bfm:reset

	soc_system soc_system_inst (
		.clk_clk                               (soc_system_inst_clk_bfm_clk_clk),                                   //                       clk.clk
		.reset_reset_n                         (soc_system_inst_reset_bfm_reset_reset),                             //                     reset.reset_n
		.memory_mem_a                          (soc_system_inst_memory_mem_a),                                      //                    memory.mem_a
		.memory_mem_ba                         (soc_system_inst_memory_mem_ba),                                     //                          .mem_ba
		.memory_mem_ck                         (soc_system_inst_memory_mem_ck),                                     //                          .mem_ck
		.memory_mem_ck_n                       (soc_system_inst_memory_mem_ck_n),                                   //                          .mem_ck_n
		.memory_mem_cke                        (soc_system_inst_memory_mem_cke),                                    //                          .mem_cke
		.memory_mem_cs_n                       (soc_system_inst_memory_mem_cs_n),                                   //                          .mem_cs_n
		.memory_mem_ras_n                      (soc_system_inst_memory_mem_ras_n),                                  //                          .mem_ras_n
		.memory_mem_cas_n                      (soc_system_inst_memory_mem_cas_n),                                  //                          .mem_cas_n
		.memory_mem_we_n                       (soc_system_inst_memory_mem_we_n),                                   //                          .mem_we_n
		.memory_mem_reset_n                    (soc_system_inst_memory_mem_reset_n),                                //                          .mem_reset_n
		.memory_mem_dq                         (soc_system_inst_memory_mem_dq),                                     //                          .mem_dq
		.memory_mem_dqs                        (soc_system_inst_memory_mem_dqs),                                    //                          .mem_dqs
		.memory_mem_dqs_n                      (soc_system_inst_memory_mem_dqs_n),                                  //                          .mem_dqs_n
		.memory_mem_odt                        (soc_system_inst_memory_mem_odt),                                    //                          .mem_odt
		.memory_mem_dm                         (soc_system_inst_memory_mem_dm),                                     //                          .mem_dm
		.memory_oct_rzqin                      (soc_system_inst_memory_bfm_conduit_oct_rzqin),                      //                          .oct_rzqin
		.hps_0_hps_io_hps_io_emac1_inst_TX_CLK (soc_system_inst_hps_0_hps_io_hps_io_emac1_inst_tx_clk),             //              hps_0_hps_io.hps_io_emac1_inst_TX_CLK
		.hps_0_hps_io_hps_io_emac1_inst_TXD0   (soc_system_inst_hps_0_hps_io_hps_io_emac1_inst_txd0),               //                          .hps_io_emac1_inst_TXD0
		.hps_0_hps_io_hps_io_emac1_inst_TXD1   (soc_system_inst_hps_0_hps_io_hps_io_emac1_inst_txd1),               //                          .hps_io_emac1_inst_TXD1
		.hps_0_hps_io_hps_io_emac1_inst_TXD2   (soc_system_inst_hps_0_hps_io_hps_io_emac1_inst_txd2),               //                          .hps_io_emac1_inst_TXD2
		.hps_0_hps_io_hps_io_emac1_inst_TXD3   (soc_system_inst_hps_0_hps_io_hps_io_emac1_inst_txd3),               //                          .hps_io_emac1_inst_TXD3
		.hps_0_hps_io_hps_io_emac1_inst_RXD0   (soc_system_inst_hps_0_hps_io_bfm_conduit_hps_io_emac1_inst_rxd0),   //                          .hps_io_emac1_inst_RXD0
		.hps_0_hps_io_hps_io_emac1_inst_MDIO   (soc_system_inst_hps_0_hps_io_hps_io_emac1_inst_mdio),               //                          .hps_io_emac1_inst_MDIO
		.hps_0_hps_io_hps_io_emac1_inst_MDC    (soc_system_inst_hps_0_hps_io_hps_io_emac1_inst_mdc),                //                          .hps_io_emac1_inst_MDC
		.hps_0_hps_io_hps_io_emac1_inst_RX_CTL (soc_system_inst_hps_0_hps_io_bfm_conduit_hps_io_emac1_inst_rx_ctl), //                          .hps_io_emac1_inst_RX_CTL
		.hps_0_hps_io_hps_io_emac1_inst_TX_CTL (soc_system_inst_hps_0_hps_io_hps_io_emac1_inst_tx_ctl),             //                          .hps_io_emac1_inst_TX_CTL
		.hps_0_hps_io_hps_io_emac1_inst_RX_CLK (soc_system_inst_hps_0_hps_io_bfm_conduit_hps_io_emac1_inst_rx_clk), //                          .hps_io_emac1_inst_RX_CLK
		.hps_0_hps_io_hps_io_emac1_inst_RXD1   (soc_system_inst_hps_0_hps_io_bfm_conduit_hps_io_emac1_inst_rxd1),   //                          .hps_io_emac1_inst_RXD1
		.hps_0_hps_io_hps_io_emac1_inst_RXD2   (soc_system_inst_hps_0_hps_io_bfm_conduit_hps_io_emac1_inst_rxd2),   //                          .hps_io_emac1_inst_RXD2
		.hps_0_hps_io_hps_io_emac1_inst_RXD3   (soc_system_inst_hps_0_hps_io_bfm_conduit_hps_io_emac1_inst_rxd3),   //                          .hps_io_emac1_inst_RXD3
		.hps_0_hps_io_hps_io_qspi_inst_IO0     (soc_system_inst_hps_0_hps_io_hps_io_qspi_inst_io0),                 //                          .hps_io_qspi_inst_IO0
		.hps_0_hps_io_hps_io_qspi_inst_IO1     (soc_system_inst_hps_0_hps_io_hps_io_qspi_inst_io1),                 //                          .hps_io_qspi_inst_IO1
		.hps_0_hps_io_hps_io_qspi_inst_IO2     (soc_system_inst_hps_0_hps_io_hps_io_qspi_inst_io2),                 //                          .hps_io_qspi_inst_IO2
		.hps_0_hps_io_hps_io_qspi_inst_IO3     (soc_system_inst_hps_0_hps_io_hps_io_qspi_inst_io3),                 //                          .hps_io_qspi_inst_IO3
		.hps_0_hps_io_hps_io_qspi_inst_SS0     (soc_system_inst_hps_0_hps_io_hps_io_qspi_inst_ss0),                 //                          .hps_io_qspi_inst_SS0
		.hps_0_hps_io_hps_io_qspi_inst_CLK     (soc_system_inst_hps_0_hps_io_hps_io_qspi_inst_clk),                 //                          .hps_io_qspi_inst_CLK
		.hps_0_hps_io_hps_io_sdio_inst_CMD     (soc_system_inst_hps_0_hps_io_hps_io_sdio_inst_cmd),                 //                          .hps_io_sdio_inst_CMD
		.hps_0_hps_io_hps_io_sdio_inst_D0      (soc_system_inst_hps_0_hps_io_hps_io_sdio_inst_d0),                  //                          .hps_io_sdio_inst_D0
		.hps_0_hps_io_hps_io_sdio_inst_D1      (soc_system_inst_hps_0_hps_io_hps_io_sdio_inst_d1),                  //                          .hps_io_sdio_inst_D1
		.hps_0_hps_io_hps_io_sdio_inst_CLK     (soc_system_inst_hps_0_hps_io_hps_io_sdio_inst_clk),                 //                          .hps_io_sdio_inst_CLK
		.hps_0_hps_io_hps_io_sdio_inst_D2      (soc_system_inst_hps_0_hps_io_hps_io_sdio_inst_d2),                  //                          .hps_io_sdio_inst_D2
		.hps_0_hps_io_hps_io_sdio_inst_D3      (soc_system_inst_hps_0_hps_io_hps_io_sdio_inst_d3),                  //                          .hps_io_sdio_inst_D3
		.hps_0_hps_io_hps_io_usb1_inst_D0      (soc_system_inst_hps_0_hps_io_hps_io_usb1_inst_d0),                  //                          .hps_io_usb1_inst_D0
		.hps_0_hps_io_hps_io_usb1_inst_D1      (soc_system_inst_hps_0_hps_io_hps_io_usb1_inst_d1),                  //                          .hps_io_usb1_inst_D1
		.hps_0_hps_io_hps_io_usb1_inst_D2      (soc_system_inst_hps_0_hps_io_hps_io_usb1_inst_d2),                  //                          .hps_io_usb1_inst_D2
		.hps_0_hps_io_hps_io_usb1_inst_D3      (soc_system_inst_hps_0_hps_io_hps_io_usb1_inst_d3),                  //                          .hps_io_usb1_inst_D3
		.hps_0_hps_io_hps_io_usb1_inst_D4      (soc_system_inst_hps_0_hps_io_hps_io_usb1_inst_d4),                  //                          .hps_io_usb1_inst_D4
		.hps_0_hps_io_hps_io_usb1_inst_D5      (soc_system_inst_hps_0_hps_io_hps_io_usb1_inst_d5),                  //                          .hps_io_usb1_inst_D5
		.hps_0_hps_io_hps_io_usb1_inst_D6      (soc_system_inst_hps_0_hps_io_hps_io_usb1_inst_d6),                  //                          .hps_io_usb1_inst_D6
		.hps_0_hps_io_hps_io_usb1_inst_D7      (soc_system_inst_hps_0_hps_io_hps_io_usb1_inst_d7),                  //                          .hps_io_usb1_inst_D7
		.hps_0_hps_io_hps_io_usb1_inst_CLK     (soc_system_inst_hps_0_hps_io_bfm_conduit_hps_io_usb1_inst_clk),     //                          .hps_io_usb1_inst_CLK
		.hps_0_hps_io_hps_io_usb1_inst_STP     (soc_system_inst_hps_0_hps_io_hps_io_usb1_inst_stp),                 //                          .hps_io_usb1_inst_STP
		.hps_0_hps_io_hps_io_usb1_inst_DIR     (soc_system_inst_hps_0_hps_io_bfm_conduit_hps_io_usb1_inst_dir),     //                          .hps_io_usb1_inst_DIR
		.hps_0_hps_io_hps_io_usb1_inst_NXT     (soc_system_inst_hps_0_hps_io_bfm_conduit_hps_io_usb1_inst_nxt),     //                          .hps_io_usb1_inst_NXT
		.hps_0_hps_io_hps_io_spim0_inst_CLK    (soc_system_inst_hps_0_hps_io_hps_io_spim0_inst_clk),                //                          .hps_io_spim0_inst_CLK
		.hps_0_hps_io_hps_io_spim0_inst_MOSI   (soc_system_inst_hps_0_hps_io_hps_io_spim0_inst_mosi),               //                          .hps_io_spim0_inst_MOSI
		.hps_0_hps_io_hps_io_spim0_inst_MISO   (soc_system_inst_hps_0_hps_io_bfm_conduit_hps_io_spim0_inst_miso),   //                          .hps_io_spim0_inst_MISO
		.hps_0_hps_io_hps_io_spim0_inst_SS0    (soc_system_inst_hps_0_hps_io_hps_io_spim0_inst_ss0),                //                          .hps_io_spim0_inst_SS0
		.hps_0_hps_io_hps_io_spim1_inst_CLK    (soc_system_inst_hps_0_hps_io_hps_io_spim1_inst_clk),                //                          .hps_io_spim1_inst_CLK
		.hps_0_hps_io_hps_io_spim1_inst_MOSI   (soc_system_inst_hps_0_hps_io_hps_io_spim1_inst_mosi),               //                          .hps_io_spim1_inst_MOSI
		.hps_0_hps_io_hps_io_spim1_inst_MISO   (soc_system_inst_hps_0_hps_io_bfm_conduit_hps_io_spim1_inst_miso),   //                          .hps_io_spim1_inst_MISO
		.hps_0_hps_io_hps_io_spim1_inst_SS0    (soc_system_inst_hps_0_hps_io_hps_io_spim1_inst_ss0),                //                          .hps_io_spim1_inst_SS0
		.hps_0_hps_io_hps_io_uart0_inst_RX     (soc_system_inst_hps_0_hps_io_bfm_conduit_hps_io_uart0_inst_rx),     //                          .hps_io_uart0_inst_RX
		.hps_0_hps_io_hps_io_uart0_inst_TX     (soc_system_inst_hps_0_hps_io_hps_io_uart0_inst_tx),                 //                          .hps_io_uart0_inst_TX
		.hps_0_hps_io_hps_io_i2c1_inst_SDA     (soc_system_inst_hps_0_hps_io_hps_io_i2c1_inst_sda),                 //                          .hps_io_i2c1_inst_SDA
		.hps_0_hps_io_hps_io_i2c1_inst_SCL     (soc_system_inst_hps_0_hps_io_hps_io_i2c1_inst_scl),                 //                          .hps_io_i2c1_inst_SCL
		.hps_0_hps_io_hps_io_gpio_inst_GPIO00  (soc_system_inst_hps_0_hps_io_hps_io_gpio_inst_gpio00),              //                          .hps_io_gpio_inst_GPIO00
		.hps_0_hps_io_hps_io_gpio_inst_GPIO09  (soc_system_inst_hps_0_hps_io_hps_io_gpio_inst_gpio09),              //                          .hps_io_gpio_inst_GPIO09
		.hps_0_hps_io_hps_io_gpio_inst_GPIO35  (soc_system_inst_hps_0_hps_io_hps_io_gpio_inst_gpio35),              //                          .hps_io_gpio_inst_GPIO35
		.hps_0_hps_io_hps_io_gpio_inst_GPIO40  (soc_system_inst_hps_0_hps_io_hps_io_gpio_inst_gpio40),              //                          .hps_io_gpio_inst_GPIO40
		.hps_0_hps_io_hps_io_gpio_inst_GPIO48  (soc_system_inst_hps_0_hps_io_hps_io_gpio_inst_gpio48),              //                          .hps_io_gpio_inst_GPIO48
		.hps_0_hps_io_hps_io_gpio_inst_GPIO53  (soc_system_inst_hps_0_hps_io_hps_io_gpio_inst_gpio53),              //                          .hps_io_gpio_inst_GPIO53
		.hps_0_hps_io_hps_io_gpio_inst_GPIO54  (soc_system_inst_hps_0_hps_io_hps_io_gpio_inst_gpio54),              //                          .hps_io_gpio_inst_GPIO54
		.hps_0_hps_io_hps_io_gpio_inst_GPIO55  (soc_system_inst_hps_0_hps_io_hps_io_gpio_inst_gpio55),              //                          .hps_io_gpio_inst_GPIO55
		.hps_0_hps_io_hps_io_gpio_inst_GPIO56  (soc_system_inst_hps_0_hps_io_hps_io_gpio_inst_gpio56),              //                          .hps_io_gpio_inst_GPIO56
		.hps_0_hps_io_hps_io_gpio_inst_GPIO61  (soc_system_inst_hps_0_hps_io_hps_io_gpio_inst_gpio61),              //                          .hps_io_gpio_inst_GPIO61
		.hps_0_hps_io_hps_io_gpio_inst_GPIO62  (soc_system_inst_hps_0_hps_io_hps_io_gpio_inst_gpio62),              //                          .hps_io_gpio_inst_GPIO62
		.hps_0_f2h_stm_hw_events_stm_hwevents  (soc_system_inst_hps_0_f2h_stm_hw_events_bfm_conduit_stm_hwevents),  //   hps_0_f2h_stm_hw_events.stm_hwevents
		.hps_0_f2h_warm_reset_req_reset_n      (soc_system_inst_hps_0_f2h_warm_reset_req_bfm_reset_reset),          //  hps_0_f2h_warm_reset_req.reset_n
		.hps_0_f2h_debug_reset_req_reset_n     (soc_system_inst_hps_0_f2h_debug_reset_req_bfm_reset_reset),         // hps_0_f2h_debug_reset_req.reset_n
		.hps_0_f2h_cold_reset_req_reset_n      (soc_system_inst_hps_0_f2h_cold_reset_req_bfm_reset_reset),          //  hps_0_f2h_cold_reset_req.reset_n
		.reg_avl_waitrequest                   (soc_system_inst_reg_avl_waitrequest),                               //                   reg_avl.waitrequest
		.reg_avl_readdata                      (soc_system_inst_reg_avl_readdata),                                  //                          .readdata
		.reg_avl_readdatavalid                 (soc_system_inst_reg_avl_readdatavalid),                             //                          .readdatavalid
		.reg_avl_burstcount                    (soc_system_inst_reg_avl_burstcount),                                //                          .burstcount
		.reg_avl_writedata                     (soc_system_inst_reg_avl_writedata),                                 //                          .writedata
		.reg_avl_address                       (soc_system_inst_reg_avl_address),                                   //                          .address
		.reg_avl_write                         (soc_system_inst_reg_avl_write),                                     //                          .write
		.reg_avl_read                          (soc_system_inst_reg_avl_read),                                      //                          .read
		.reg_avl_byteenable                    (soc_system_inst_reg_avl_byteenable),                                //                          .byteenable
		.reg_avl_debugaccess                   (soc_system_inst_reg_avl_debugaccess),                               //                          .debugaccess
		.hps_0_h2f_reset_reset_n               (),                                                                  //           hps_0_h2f_reset.reset_n
		.h2f_0_waitrequest                     (soc_system_inst_h2f_0_waitrequest),                                 //                     h2f_0.waitrequest
		.h2f_0_readdata                        (soc_system_inst_h2f_0_readdata),                                    //                          .readdata
		.h2f_0_readdatavalid                   (soc_system_inst_h2f_0_readdatavalid),                               //                          .readdatavalid
		.h2f_0_burstcount                      (soc_system_inst_h2f_0_burstcount),                                  //                          .burstcount
		.h2f_0_writedata                       (soc_system_inst_h2f_0_writedata),                                   //                          .writedata
		.h2f_0_address                         (soc_system_inst_h2f_0_address),                                     //                          .address
		.h2f_0_write                           (soc_system_inst_h2f_0_write),                                       //                          .write
		.h2f_0_read                            (soc_system_inst_h2f_0_read),                                        //                          .read
		.h2f_0_byteenable                      (soc_system_inst_h2f_0_byteenable),                                  //                          .byteenable
		.h2f_0_debugaccess                     (soc_system_inst_h2f_0_debugaccess),                                 //                          .debugaccess
		.afi_clk_clk                           (soc_system_inst_afi_clk_bfm_clk_clk)                                //                   afi_clk.clk
	);

	altera_avalon_clock_source #(
		.CLOCK_RATE (50000000),
		.CLOCK_UNIT (1)
	) soc_system_inst_clk_bfm (
		.clk (soc_system_inst_clk_bfm_clk_clk)  // clk.clk
	);

	altera_avalon_clock_source #(
		.CLOCK_RATE (50000000),
		.CLOCK_UNIT (1)
	) soc_system_inst_afi_clk_bfm (
		.clk (soc_system_inst_afi_clk_bfm_clk_clk)  // clk.clk
	);

	altera_avalon_reset_source #(
		.ASSERT_HIGH_RESET    (0),
		.INITIAL_RESET_CYCLES (50)
	) soc_system_inst_reset_bfm (
		.reset (soc_system_inst_reset_bfm_reset_reset), // reset.reset_n
		.clk   (soc_system_inst_clk_bfm_clk_clk)        //   clk.clk
	);

	altera_avalon_reset_source #(
		.ASSERT_HIGH_RESET    (0),
		.INITIAL_RESET_CYCLES (50)
	) soc_system_inst_hps_0_f2h_warm_reset_req_bfm (
		.reset (soc_system_inst_hps_0_f2h_warm_reset_req_bfm_reset_reset), // reset.reset_n
		.clk   (soc_system_inst_clk_bfm_clk_clk)                           //   clk.clk
	);

	altera_avalon_reset_source #(
		.ASSERT_HIGH_RESET    (0),
		.INITIAL_RESET_CYCLES (50)
	) soc_system_inst_hps_0_f2h_debug_reset_req_bfm (
		.reset (soc_system_inst_hps_0_f2h_debug_reset_req_bfm_reset_reset), // reset.reset_n
		.clk   (soc_system_inst_clk_bfm_clk_clk)                            //   clk.clk
	);

	altera_avalon_reset_source #(
		.ASSERT_HIGH_RESET    (0),
		.INITIAL_RESET_CYCLES (50)
	) soc_system_inst_hps_0_f2h_cold_reset_req_bfm (
		.reset (soc_system_inst_hps_0_f2h_cold_reset_req_bfm_reset_reset), // reset.reset_n
		.clk   (soc_system_inst_clk_bfm_clk_clk)                           //   clk.clk
	);

	altera_conduit_bfm soc_system_inst_memory_bfm (
		.sig_mem_a       (soc_system_inst_memory_mem_a),                 // conduit.mem_a
		.sig_mem_ba      (soc_system_inst_memory_mem_ba),                //        .mem_ba
		.sig_mem_ck      (soc_system_inst_memory_mem_ck),                //        .mem_ck
		.sig_mem_ck_n    (soc_system_inst_memory_mem_ck_n),              //        .mem_ck_n
		.sig_mem_cke     (soc_system_inst_memory_mem_cke),               //        .mem_cke
		.sig_mem_cs_n    (soc_system_inst_memory_mem_cs_n),              //        .mem_cs_n
		.sig_mem_ras_n   (soc_system_inst_memory_mem_ras_n),             //        .mem_ras_n
		.sig_mem_cas_n   (soc_system_inst_memory_mem_cas_n),             //        .mem_cas_n
		.sig_mem_we_n    (soc_system_inst_memory_mem_we_n),              //        .mem_we_n
		.sig_mem_reset_n (soc_system_inst_memory_mem_reset_n),           //        .mem_reset_n
		.sig_mem_dq      (soc_system_inst_memory_mem_dq),                //        .mem_dq
		.sig_mem_dqs     (soc_system_inst_memory_mem_dqs),               //        .mem_dqs
		.sig_mem_dqs_n   (soc_system_inst_memory_mem_dqs_n),             //        .mem_dqs_n
		.sig_mem_odt     (soc_system_inst_memory_mem_odt),               //        .mem_odt
		.sig_mem_dm      (soc_system_inst_memory_mem_dm),                //        .mem_dm
		.sig_oct_rzqin   (soc_system_inst_memory_bfm_conduit_oct_rzqin)  //        .oct_rzqin
	);

	altera_conduit_bfm_0002 soc_system_inst_hps_0_hps_io_bfm (
		.sig_hps_io_emac1_inst_TX_CLK (soc_system_inst_hps_0_hps_io_hps_io_emac1_inst_tx_clk),             // conduit.hps_io_emac1_inst_TX_CLK
		.sig_hps_io_emac1_inst_TXD0   (soc_system_inst_hps_0_hps_io_hps_io_emac1_inst_txd0),               //        .hps_io_emac1_inst_TXD0
		.sig_hps_io_emac1_inst_TXD1   (soc_system_inst_hps_0_hps_io_hps_io_emac1_inst_txd1),               //        .hps_io_emac1_inst_TXD1
		.sig_hps_io_emac1_inst_TXD2   (soc_system_inst_hps_0_hps_io_hps_io_emac1_inst_txd2),               //        .hps_io_emac1_inst_TXD2
		.sig_hps_io_emac1_inst_TXD3   (soc_system_inst_hps_0_hps_io_hps_io_emac1_inst_txd3),               //        .hps_io_emac1_inst_TXD3
		.sig_hps_io_emac1_inst_RXD0   (soc_system_inst_hps_0_hps_io_bfm_conduit_hps_io_emac1_inst_rxd0),   //        .hps_io_emac1_inst_RXD0
		.sig_hps_io_emac1_inst_MDIO   (soc_system_inst_hps_0_hps_io_hps_io_emac1_inst_mdio),               //        .hps_io_emac1_inst_MDIO
		.sig_hps_io_emac1_inst_MDC    (soc_system_inst_hps_0_hps_io_hps_io_emac1_inst_mdc),                //        .hps_io_emac1_inst_MDC
		.sig_hps_io_emac1_inst_RX_CTL (soc_system_inst_hps_0_hps_io_bfm_conduit_hps_io_emac1_inst_rx_ctl), //        .hps_io_emac1_inst_RX_CTL
		.sig_hps_io_emac1_inst_TX_CTL (soc_system_inst_hps_0_hps_io_hps_io_emac1_inst_tx_ctl),             //        .hps_io_emac1_inst_TX_CTL
		.sig_hps_io_emac1_inst_RX_CLK (soc_system_inst_hps_0_hps_io_bfm_conduit_hps_io_emac1_inst_rx_clk), //        .hps_io_emac1_inst_RX_CLK
		.sig_hps_io_emac1_inst_RXD1   (soc_system_inst_hps_0_hps_io_bfm_conduit_hps_io_emac1_inst_rxd1),   //        .hps_io_emac1_inst_RXD1
		.sig_hps_io_emac1_inst_RXD2   (soc_system_inst_hps_0_hps_io_bfm_conduit_hps_io_emac1_inst_rxd2),   //        .hps_io_emac1_inst_RXD2
		.sig_hps_io_emac1_inst_RXD3   (soc_system_inst_hps_0_hps_io_bfm_conduit_hps_io_emac1_inst_rxd3),   //        .hps_io_emac1_inst_RXD3
		.sig_hps_io_qspi_inst_IO0     (soc_system_inst_hps_0_hps_io_hps_io_qspi_inst_io0),                 //        .hps_io_qspi_inst_IO0
		.sig_hps_io_qspi_inst_IO1     (soc_system_inst_hps_0_hps_io_hps_io_qspi_inst_io1),                 //        .hps_io_qspi_inst_IO1
		.sig_hps_io_qspi_inst_IO2     (soc_system_inst_hps_0_hps_io_hps_io_qspi_inst_io2),                 //        .hps_io_qspi_inst_IO2
		.sig_hps_io_qspi_inst_IO3     (soc_system_inst_hps_0_hps_io_hps_io_qspi_inst_io3),                 //        .hps_io_qspi_inst_IO3
		.sig_hps_io_qspi_inst_SS0     (soc_system_inst_hps_0_hps_io_hps_io_qspi_inst_ss0),                 //        .hps_io_qspi_inst_SS0
		.sig_hps_io_qspi_inst_CLK     (soc_system_inst_hps_0_hps_io_hps_io_qspi_inst_clk),                 //        .hps_io_qspi_inst_CLK
		.sig_hps_io_sdio_inst_CMD     (soc_system_inst_hps_0_hps_io_hps_io_sdio_inst_cmd),                 //        .hps_io_sdio_inst_CMD
		.sig_hps_io_sdio_inst_D0      (soc_system_inst_hps_0_hps_io_hps_io_sdio_inst_d0),                  //        .hps_io_sdio_inst_D0
		.sig_hps_io_sdio_inst_D1      (soc_system_inst_hps_0_hps_io_hps_io_sdio_inst_d1),                  //        .hps_io_sdio_inst_D1
		.sig_hps_io_sdio_inst_CLK     (soc_system_inst_hps_0_hps_io_hps_io_sdio_inst_clk),                 //        .hps_io_sdio_inst_CLK
		.sig_hps_io_sdio_inst_D2      (soc_system_inst_hps_0_hps_io_hps_io_sdio_inst_d2),                  //        .hps_io_sdio_inst_D2
		.sig_hps_io_sdio_inst_D3      (soc_system_inst_hps_0_hps_io_hps_io_sdio_inst_d3),                  //        .hps_io_sdio_inst_D3
		.sig_hps_io_usb1_inst_D0      (soc_system_inst_hps_0_hps_io_hps_io_usb1_inst_d0),                  //        .hps_io_usb1_inst_D0
		.sig_hps_io_usb1_inst_D1      (soc_system_inst_hps_0_hps_io_hps_io_usb1_inst_d1),                  //        .hps_io_usb1_inst_D1
		.sig_hps_io_usb1_inst_D2      (soc_system_inst_hps_0_hps_io_hps_io_usb1_inst_d2),                  //        .hps_io_usb1_inst_D2
		.sig_hps_io_usb1_inst_D3      (soc_system_inst_hps_0_hps_io_hps_io_usb1_inst_d3),                  //        .hps_io_usb1_inst_D3
		.sig_hps_io_usb1_inst_D4      (soc_system_inst_hps_0_hps_io_hps_io_usb1_inst_d4),                  //        .hps_io_usb1_inst_D4
		.sig_hps_io_usb1_inst_D5      (soc_system_inst_hps_0_hps_io_hps_io_usb1_inst_d5),                  //        .hps_io_usb1_inst_D5
		.sig_hps_io_usb1_inst_D6      (soc_system_inst_hps_0_hps_io_hps_io_usb1_inst_d6),                  //        .hps_io_usb1_inst_D6
		.sig_hps_io_usb1_inst_D7      (soc_system_inst_hps_0_hps_io_hps_io_usb1_inst_d7),                  //        .hps_io_usb1_inst_D7
		.sig_hps_io_usb1_inst_CLK     (soc_system_inst_hps_0_hps_io_bfm_conduit_hps_io_usb1_inst_clk),     //        .hps_io_usb1_inst_CLK
		.sig_hps_io_usb1_inst_STP     (soc_system_inst_hps_0_hps_io_hps_io_usb1_inst_stp),                 //        .hps_io_usb1_inst_STP
		.sig_hps_io_usb1_inst_DIR     (soc_system_inst_hps_0_hps_io_bfm_conduit_hps_io_usb1_inst_dir),     //        .hps_io_usb1_inst_DIR
		.sig_hps_io_usb1_inst_NXT     (soc_system_inst_hps_0_hps_io_bfm_conduit_hps_io_usb1_inst_nxt),     //        .hps_io_usb1_inst_NXT
		.sig_hps_io_spim0_inst_CLK    (soc_system_inst_hps_0_hps_io_hps_io_spim0_inst_clk),                //        .hps_io_spim0_inst_CLK
		.sig_hps_io_spim0_inst_MOSI   (soc_system_inst_hps_0_hps_io_hps_io_spim0_inst_mosi),               //        .hps_io_spim0_inst_MOSI
		.sig_hps_io_spim0_inst_MISO   (soc_system_inst_hps_0_hps_io_bfm_conduit_hps_io_spim0_inst_miso),   //        .hps_io_spim0_inst_MISO
		.sig_hps_io_spim0_inst_SS0    (soc_system_inst_hps_0_hps_io_hps_io_spim0_inst_ss0),                //        .hps_io_spim0_inst_SS0
		.sig_hps_io_spim1_inst_CLK    (soc_system_inst_hps_0_hps_io_hps_io_spim1_inst_clk),                //        .hps_io_spim1_inst_CLK
		.sig_hps_io_spim1_inst_MOSI   (soc_system_inst_hps_0_hps_io_hps_io_spim1_inst_mosi),               //        .hps_io_spim1_inst_MOSI
		.sig_hps_io_spim1_inst_MISO   (soc_system_inst_hps_0_hps_io_bfm_conduit_hps_io_spim1_inst_miso),   //        .hps_io_spim1_inst_MISO
		.sig_hps_io_spim1_inst_SS0    (soc_system_inst_hps_0_hps_io_hps_io_spim1_inst_ss0),                //        .hps_io_spim1_inst_SS0
		.sig_hps_io_uart0_inst_RX     (soc_system_inst_hps_0_hps_io_bfm_conduit_hps_io_uart0_inst_rx),     //        .hps_io_uart0_inst_RX
		.sig_hps_io_uart0_inst_TX     (soc_system_inst_hps_0_hps_io_hps_io_uart0_inst_tx),                 //        .hps_io_uart0_inst_TX
		.sig_hps_io_i2c1_inst_SDA     (soc_system_inst_hps_0_hps_io_hps_io_i2c1_inst_sda),                 //        .hps_io_i2c1_inst_SDA
		.sig_hps_io_i2c1_inst_SCL     (soc_system_inst_hps_0_hps_io_hps_io_i2c1_inst_scl),                 //        .hps_io_i2c1_inst_SCL
		.sig_hps_io_gpio_inst_GPIO00  (soc_system_inst_hps_0_hps_io_hps_io_gpio_inst_gpio00),              //        .hps_io_gpio_inst_GPIO00
		.sig_hps_io_gpio_inst_GPIO09  (soc_system_inst_hps_0_hps_io_hps_io_gpio_inst_gpio09),              //        .hps_io_gpio_inst_GPIO09
		.sig_hps_io_gpio_inst_GPIO35  (soc_system_inst_hps_0_hps_io_hps_io_gpio_inst_gpio35),              //        .hps_io_gpio_inst_GPIO35
		.sig_hps_io_gpio_inst_GPIO40  (soc_system_inst_hps_0_hps_io_hps_io_gpio_inst_gpio40),              //        .hps_io_gpio_inst_GPIO40
		.sig_hps_io_gpio_inst_GPIO48  (soc_system_inst_hps_0_hps_io_hps_io_gpio_inst_gpio48),              //        .hps_io_gpio_inst_GPIO48
		.sig_hps_io_gpio_inst_GPIO53  (soc_system_inst_hps_0_hps_io_hps_io_gpio_inst_gpio53),              //        .hps_io_gpio_inst_GPIO53
		.sig_hps_io_gpio_inst_GPIO54  (soc_system_inst_hps_0_hps_io_hps_io_gpio_inst_gpio54),              //        .hps_io_gpio_inst_GPIO54
		.sig_hps_io_gpio_inst_GPIO55  (soc_system_inst_hps_0_hps_io_hps_io_gpio_inst_gpio55),              //        .hps_io_gpio_inst_GPIO55
		.sig_hps_io_gpio_inst_GPIO56  (soc_system_inst_hps_0_hps_io_hps_io_gpio_inst_gpio56),              //        .hps_io_gpio_inst_GPIO56
		.sig_hps_io_gpio_inst_GPIO61  (soc_system_inst_hps_0_hps_io_hps_io_gpio_inst_gpio61),              //        .hps_io_gpio_inst_GPIO61
		.sig_hps_io_gpio_inst_GPIO62  (soc_system_inst_hps_0_hps_io_hps_io_gpio_inst_gpio62)               //        .hps_io_gpio_inst_GPIO62
	);

	altera_conduit_bfm_0003 soc_system_inst_hps_0_f2h_stm_hw_events_bfm (
		.sig_stm_hwevents (soc_system_inst_hps_0_f2h_stm_hw_events_bfm_conduit_stm_hwevents)  // conduit.stm_hwevents
	);

	altera_avalon_mm_slave_bfm #(
		.AV_ADDRESS_W               (10),
		.AV_SYMBOL_W                (8),
		.AV_NUMSYMBOLS              (4),
		.AV_BURSTCOUNT_W            (1),
		.AV_READRESPONSE_W          (1),
		.AV_WRITERESPONSE_W         (1),
		.USE_READ                   (1),
		.USE_WRITE                  (1),
		.USE_ADDRESS                (1),
		.USE_BYTE_ENABLE            (1),
		.USE_BURSTCOUNT             (1),
		.USE_READ_DATA              (1),
		.USE_READ_DATA_VALID        (1),
		.USE_WRITE_DATA             (1),
		.USE_BEGIN_TRANSFER         (0),
		.USE_BEGIN_BURST_TRANSFER   (0),
		.USE_WAIT_REQUEST           (1),
		.USE_TRANSACTIONID          (0),
		.USE_WRITERESPONSE          (0),
		.USE_READRESPONSE           (0),
		.USE_CLKEN                  (0),
		.AV_BURST_LINEWRAP          (0),
		.AV_BURST_BNDR_ONLY         (0),
		.AV_MAX_PENDING_READS       (64),
		.AV_MAX_PENDING_WRITES      (0),
		.AV_FIX_READ_LATENCY        (0),
		.AV_READ_WAIT_TIME          (1),
		.AV_WRITE_WAIT_TIME         (0),
		.REGISTER_WAITREQUEST       (0),
		.AV_REGISTERINCOMINGSIGNALS (0),
		.VHDL_ID                    (0)
	) soc_system_inst_reg_avl_bfm (
		.clk                      (soc_system_inst_clk_bfm_clk_clk),        //       clk.clk
		.reset                    (~soc_system_inst_reset_bfm_reset_reset), // clk_reset.reset
		.avs_writedata            (soc_system_inst_reg_avl_writedata),      //        s0.writedata
		.avs_burstcount           (soc_system_inst_reg_avl_burstcount),     //          .burstcount
		.avs_readdata             (soc_system_inst_reg_avl_readdata),       //          .readdata
		.avs_address              (soc_system_inst_reg_avl_address),        //          .address
		.avs_waitrequest          (soc_system_inst_reg_avl_waitrequest),    //          .waitrequest
		.avs_write                (soc_system_inst_reg_avl_write),          //          .write
		.avs_read                 (soc_system_inst_reg_avl_read),           //          .read
		.avs_byteenable           (soc_system_inst_reg_avl_byteenable),     //          .byteenable
		.avs_readdatavalid        (soc_system_inst_reg_avl_readdatavalid),  //          .readdatavalid
		.avs_debugaccess          (soc_system_inst_reg_avl_debugaccess),    //          .debugaccess
		.avs_begintransfer        (1'b0),                                   // (terminated)
		.avs_beginbursttransfer   (1'b0),                                   // (terminated)
		.avs_arbiterlock          (1'b0),                                   // (terminated)
		.avs_lock                 (1'b0),                                   // (terminated)
		.avs_transactionid        (8'b00000000),                            // (terminated)
		.avs_readid               (),                                       // (terminated)
		.avs_writeid              (),                                       // (terminated)
		.avs_clken                (1'b1),                                   // (terminated)
		.avs_response             (),                                       // (terminated)
		.avs_writeresponserequest (1'b0),                                   // (terminated)
		.avs_writeresponsevalid   (),                                       // (terminated)
		.avs_readresponse         (),                                       // (terminated)
		.avs_writeresponse        ()                                        // (terminated)
	);

	altera_avalon_mm_slave_bfm #(
		.AV_ADDRESS_W               (26),
		.AV_SYMBOL_W                (8),
		.AV_NUMSYMBOLS              (16),
		.AV_BURSTCOUNT_W            (6),
		.AV_READRESPONSE_W          (1),
		.AV_WRITERESPONSE_W         (1),
		.USE_READ                   (1),
		.USE_WRITE                  (1),
		.USE_ADDRESS                (1),
		.USE_BYTE_ENABLE            (1),
		.USE_BURSTCOUNT             (1),
		.USE_READ_DATA              (1),
		.USE_READ_DATA_VALID        (1),
		.USE_WRITE_DATA             (1),
		.USE_BEGIN_TRANSFER         (0),
		.USE_BEGIN_BURST_TRANSFER   (0),
		.USE_WAIT_REQUEST           (1),
		.USE_TRANSACTIONID          (0),
		.USE_WRITERESPONSE          (0),
		.USE_READRESPONSE           (0),
		.USE_CLKEN                  (0),
		.AV_BURST_LINEWRAP          (0),
		.AV_BURST_BNDR_ONLY         (0),
		.AV_MAX_PENDING_READS       (64),
		.AV_MAX_PENDING_WRITES      (0),
		.AV_FIX_READ_LATENCY        (0),
		.AV_READ_WAIT_TIME          (1),
		.AV_WRITE_WAIT_TIME         (0),
		.REGISTER_WAITREQUEST       (0),
		.AV_REGISTERINCOMINGSIGNALS (0),
		.VHDL_ID                    (1)
	) soc_system_inst_h2f_0_bfm (
		.clk                      (soc_system_inst_afi_clk_bfm_clk_clk), //       clk.clk
		.reset                    (rst_controller_reset_out_reset),      // clk_reset.reset
		.avs_writedata            (soc_system_inst_h2f_0_writedata),     //        s0.writedata
		.avs_burstcount           (soc_system_inst_h2f_0_burstcount),    //          .burstcount
		.avs_readdata             (soc_system_inst_h2f_0_readdata),      //          .readdata
		.avs_address              (soc_system_inst_h2f_0_address),       //          .address
		.avs_waitrequest          (soc_system_inst_h2f_0_waitrequest),   //          .waitrequest
		.avs_write                (soc_system_inst_h2f_0_write),         //          .write
		.avs_read                 (soc_system_inst_h2f_0_read),          //          .read
		.avs_byteenable           (soc_system_inst_h2f_0_byteenable),    //          .byteenable
		.avs_readdatavalid        (soc_system_inst_h2f_0_readdatavalid), //          .readdatavalid
		.avs_debugaccess          (soc_system_inst_h2f_0_debugaccess),   //          .debugaccess
		.avs_begintransfer        (1'b0),                                // (terminated)
		.avs_beginbursttransfer   (1'b0),                                // (terminated)
		.avs_arbiterlock          (1'b0),                                // (terminated)
		.avs_lock                 (1'b0),                                // (terminated)
		.avs_transactionid        (8'b00000000),                         // (terminated)
		.avs_readid               (),                                    // (terminated)
		.avs_writeid              (),                                    // (terminated)
		.avs_clken                (1'b1),                                // (terminated)
		.avs_response             (),                                    // (terminated)
		.avs_writeresponserequest (1'b0),                                // (terminated)
		.avs_writeresponsevalid   (),                                    // (terminated)
		.avs_readresponse         (),                                    // (terminated)
		.avs_writeresponse        ()                                     // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~soc_system_inst_reset_bfm_reset_reset), // reset_in0.reset
		.clk            (soc_system_inst_afi_clk_bfm_clk_clk),    //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),         // reset_out.reset
		.reset_req      (),                                       // (terminated)
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_in1      (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

endmodule
